magic
tech sky130A
magscale 1 2
timestamp 1611412735
<< obsli1 >>
rect 38 31 231786 295457
<< obsm1 >>
rect 38 0 231786 295772
<< metal2 >>
rect 332 297072 388 297872
rect 3184 297072 3240 297872
rect 6128 297072 6184 297872
rect 9072 297072 9128 297872
rect 12016 297072 12072 297872
rect 14868 297072 14924 297872
rect 17812 297072 17868 297872
rect 20756 297072 20812 297872
rect 23700 297072 23756 297872
rect 26644 297072 26700 297872
rect 29496 297072 29552 297872
rect 32440 297072 32496 297872
rect 35384 297072 35440 297872
rect 38328 297072 38384 297872
rect 41272 297072 41328 297872
rect 44124 297072 44180 297872
rect 47068 297072 47124 297872
rect 50012 297072 50068 297872
rect 52956 297072 53012 297872
rect 55808 297072 55864 297872
rect 58752 297072 58808 297872
rect 61696 297072 61752 297872
rect 64640 297072 64696 297872
rect 67584 297072 67640 297872
rect 70436 297072 70492 297872
rect 73380 297072 73436 297872
rect 76324 297072 76380 297872
rect 79268 297072 79324 297872
rect 82212 297072 82268 297872
rect 85064 297072 85120 297872
rect 88008 297072 88064 297872
rect 90952 297072 91008 297872
rect 93896 297072 93952 297872
rect 96748 297072 96804 297872
rect 99692 297072 99748 297872
rect 102636 297072 102692 297872
rect 105580 297072 105636 297872
rect 108524 297072 108580 297872
rect 111376 297072 111432 297872
rect 114320 297072 114376 297872
rect 117264 297072 117320 297872
rect 120208 297072 120264 297872
rect 123152 297072 123208 297872
rect 126004 297072 126060 297872
rect 128948 297072 129004 297872
rect 131892 297072 131948 297872
rect 134836 297072 134892 297872
rect 137780 297072 137836 297872
rect 140632 297072 140688 297872
rect 143576 297072 143632 297872
rect 146520 297072 146576 297872
rect 149464 297072 149520 297872
rect 152316 297072 152372 297872
rect 155260 297072 155316 297872
rect 158204 297072 158260 297872
rect 161148 297072 161204 297872
rect 164092 297072 164148 297872
rect 166944 297072 167000 297872
rect 169888 297072 169944 297872
rect 172832 297072 172888 297872
rect 175776 297072 175832 297872
rect 178720 297072 178776 297872
rect 181572 297072 181628 297872
rect 184516 297072 184572 297872
rect 187460 297072 187516 297872
rect 190404 297072 190460 297872
rect 193256 297072 193312 297872
rect 196200 297072 196256 297872
rect 199144 297072 199200 297872
rect 202088 297072 202144 297872
rect 205032 297072 205088 297872
rect 207884 297072 207940 297872
rect 210828 297072 210884 297872
rect 213772 297072 213828 297872
rect 216716 297072 216772 297872
rect 219660 297072 219716 297872
rect 222512 297072 222568 297872
rect 225456 297072 225512 297872
rect 228400 297072 228456 297872
rect 231344 297072 231400 297872
<< obsm2 >>
rect 444 297016 3128 297072
rect 3296 297016 6072 297072
rect 6240 297016 9016 297072
rect 9184 297016 11960 297072
rect 12128 297016 14812 297072
rect 14980 297016 17756 297072
rect 17924 297016 20700 297072
rect 20868 297016 23644 297072
rect 23812 297016 26588 297072
rect 26756 297016 29440 297072
rect 29608 297016 32384 297072
rect 32552 297016 35328 297072
rect 35496 297016 38272 297072
rect 38440 297016 41216 297072
rect 41384 297016 44068 297072
rect 44236 297016 47012 297072
rect 47180 297016 49956 297072
rect 50124 297016 52900 297072
rect 53068 297016 55752 297072
rect 55920 297016 58696 297072
rect 58864 297016 61640 297072
rect 61808 297016 64584 297072
rect 64752 297016 67528 297072
rect 67696 297016 70380 297072
rect 70548 297016 73324 297072
rect 73492 297016 76268 297072
rect 76436 297016 79212 297072
rect 79380 297016 82156 297072
rect 82324 297016 85008 297072
rect 85176 297016 87952 297072
rect 88120 297016 90896 297072
rect 91064 297016 93840 297072
rect 94008 297016 96692 297072
rect 96860 297016 99636 297072
rect 99804 297016 102580 297072
rect 102748 297016 105524 297072
rect 105692 297016 108468 297072
rect 108636 297016 111320 297072
rect 111488 297016 114264 297072
rect 114432 297016 117208 297072
rect 117376 297016 120152 297072
rect 120320 297016 123096 297072
rect 123264 297016 125948 297072
rect 126116 297016 128892 297072
rect 129060 297016 131836 297072
rect 132004 297016 134780 297072
rect 134948 297016 137724 297072
rect 137892 297016 140576 297072
rect 140744 297016 143520 297072
rect 143688 297016 146464 297072
rect 146632 297016 149408 297072
rect 149576 297016 152260 297072
rect 152428 297016 155204 297072
rect 155372 297016 158148 297072
rect 158316 297016 161092 297072
rect 161260 297016 164036 297072
rect 164204 297016 166888 297072
rect 167056 297016 169832 297072
rect 170000 297016 172776 297072
rect 172944 297016 175720 297072
rect 175888 297016 178664 297072
rect 178832 297016 181516 297072
rect 181684 297016 184460 297072
rect 184628 297016 187404 297072
rect 187572 297016 190348 297072
rect 190516 297016 193200 297072
rect 193368 297016 196144 297072
rect 196312 297016 199088 297072
rect 199256 297016 202032 297072
rect 202200 297016 204976 297072
rect 205144 297016 207828 297072
rect 207996 297016 210772 297072
rect 210940 297016 213716 297072
rect 213884 297016 216660 297072
rect 216828 297016 219604 297072
rect 219772 297016 222456 297072
rect 222624 297016 225400 297072
rect 225568 297016 228344 297072
rect 228512 297016 231288 297072
rect 231456 297016 231582 297072
rect 334 0 231582 297016
<< obsm3 >>
rect 603 15 231462 295473
<< metal4 >>
rect 3142 0 3462 295488
rect 15142 0 15462 295488
rect 27142 0 27462 295488
rect 39142 0 39462 295488
rect 51142 0 51462 295488
rect 63142 0 63462 295488
rect 75142 0 75462 295488
rect 87142 0 87462 295488
rect 99142 0 99462 295488
rect 111142 0 111462 295488
rect 123142 0 123462 295488
rect 135142 0 135462 295488
rect 147142 0 147462 295488
rect 159142 0 159462 295488
rect 171142 0 171462 295488
rect 183142 0 183462 295488
rect 195142 0 195462 295488
rect 207142 0 207462 295488
rect 219142 0 219462 295488
rect 231142 0 231462 295488
<< obsm4 >>
rect 4145 8515 15062 294997
rect 15542 8515 27062 294997
rect 27542 8515 39062 294997
rect 39542 8515 51062 294997
rect 51542 8515 63062 294997
rect 63542 8515 75062 294997
rect 75542 8515 87062 294997
rect 87542 8515 99062 294997
rect 99542 8515 111062 294997
rect 111542 8515 123062 294997
rect 123542 8515 135062 294997
rect 135542 8515 147062 294997
rect 147542 8515 159062 294997
rect 159542 8515 171062 294997
rect 171542 8515 183062 294997
rect 183542 8515 195062 294997
rect 195542 8515 207062 294997
rect 207542 8515 219062 294997
rect 219542 8515 228139 294997
<< labels >>
rlabel metal2 s 93896 297072 93952 297872 6 A[0]
port 1 nsew signal input
rlabel metal2 s 96748 297072 96804 297872 6 A[1]
port 2 nsew signal input
rlabel metal2 s 99692 297072 99748 297872 6 A[2]
port 3 nsew signal input
rlabel metal2 s 102636 297072 102692 297872 6 A[3]
port 4 nsew signal input
rlabel metal2 s 105580 297072 105636 297872 6 A[4]
port 5 nsew signal input
rlabel metal2 s 108524 297072 108580 297872 6 A[5]
port 6 nsew signal input
rlabel metal2 s 111376 297072 111432 297872 6 A[6]
port 7 nsew signal input
rlabel metal2 s 114320 297072 114376 297872 6 A[7]
port 8 nsew signal input
rlabel metal2 s 117264 297072 117320 297872 6 A[8]
port 9 nsew signal input
rlabel metal2 s 120208 297072 120264 297872 6 A[9]
port 10 nsew signal input
rlabel metal2 s 123152 297072 123208 297872 6 CLK
port 11 nsew signal input
rlabel metal2 s 140632 297072 140688 297872 6 Di[0]
port 12 nsew signal input
rlabel metal2 s 169888 297072 169944 297872 6 Di[10]
port 13 nsew signal input
rlabel metal2 s 172832 297072 172888 297872 6 Di[11]
port 14 nsew signal input
rlabel metal2 s 175776 297072 175832 297872 6 Di[12]
port 15 nsew signal input
rlabel metal2 s 178720 297072 178776 297872 6 Di[13]
port 16 nsew signal input
rlabel metal2 s 181572 297072 181628 297872 6 Di[14]
port 17 nsew signal input
rlabel metal2 s 184516 297072 184572 297872 6 Di[15]
port 18 nsew signal input
rlabel metal2 s 187460 297072 187516 297872 6 Di[16]
port 19 nsew signal input
rlabel metal2 s 190404 297072 190460 297872 6 Di[17]
port 20 nsew signal input
rlabel metal2 s 193256 297072 193312 297872 6 Di[18]
port 21 nsew signal input
rlabel metal2 s 196200 297072 196256 297872 6 Di[19]
port 22 nsew signal input
rlabel metal2 s 143576 297072 143632 297872 6 Di[1]
port 23 nsew signal input
rlabel metal2 s 199144 297072 199200 297872 6 Di[20]
port 24 nsew signal input
rlabel metal2 s 202088 297072 202144 297872 6 Di[21]
port 25 nsew signal input
rlabel metal2 s 205032 297072 205088 297872 6 Di[22]
port 26 nsew signal input
rlabel metal2 s 207884 297072 207940 297872 6 Di[23]
port 27 nsew signal input
rlabel metal2 s 210828 297072 210884 297872 6 Di[24]
port 28 nsew signal input
rlabel metal2 s 213772 297072 213828 297872 6 Di[25]
port 29 nsew signal input
rlabel metal2 s 216716 297072 216772 297872 6 Di[26]
port 30 nsew signal input
rlabel metal2 s 219660 297072 219716 297872 6 Di[27]
port 31 nsew signal input
rlabel metal2 s 222512 297072 222568 297872 6 Di[28]
port 32 nsew signal input
rlabel metal2 s 225456 297072 225512 297872 6 Di[29]
port 33 nsew signal input
rlabel metal2 s 146520 297072 146576 297872 6 Di[2]
port 34 nsew signal input
rlabel metal2 s 228400 297072 228456 297872 6 Di[30]
port 35 nsew signal input
rlabel metal2 s 231344 297072 231400 297872 6 Di[31]
port 36 nsew signal input
rlabel metal2 s 149464 297072 149520 297872 6 Di[3]
port 37 nsew signal input
rlabel metal2 s 152316 297072 152372 297872 6 Di[4]
port 38 nsew signal input
rlabel metal2 s 155260 297072 155316 297872 6 Di[5]
port 39 nsew signal input
rlabel metal2 s 158204 297072 158260 297872 6 Di[6]
port 40 nsew signal input
rlabel metal2 s 161148 297072 161204 297872 6 Di[7]
port 41 nsew signal input
rlabel metal2 s 164092 297072 164148 297872 6 Di[8]
port 42 nsew signal input
rlabel metal2 s 166944 297072 167000 297872 6 Di[9]
port 43 nsew signal input
rlabel metal2 s 332 297072 388 297872 6 Do[0]
port 44 nsew signal output
rlabel metal2 s 29496 297072 29552 297872 6 Do[10]
port 45 nsew signal output
rlabel metal2 s 32440 297072 32496 297872 6 Do[11]
port 46 nsew signal output
rlabel metal2 s 35384 297072 35440 297872 6 Do[12]
port 47 nsew signal output
rlabel metal2 s 38328 297072 38384 297872 6 Do[13]
port 48 nsew signal output
rlabel metal2 s 41272 297072 41328 297872 6 Do[14]
port 49 nsew signal output
rlabel metal2 s 44124 297072 44180 297872 6 Do[15]
port 50 nsew signal output
rlabel metal2 s 47068 297072 47124 297872 6 Do[16]
port 51 nsew signal output
rlabel metal2 s 50012 297072 50068 297872 6 Do[17]
port 52 nsew signal output
rlabel metal2 s 52956 297072 53012 297872 6 Do[18]
port 53 nsew signal output
rlabel metal2 s 55808 297072 55864 297872 6 Do[19]
port 54 nsew signal output
rlabel metal2 s 3184 297072 3240 297872 6 Do[1]
port 55 nsew signal output
rlabel metal2 s 58752 297072 58808 297872 6 Do[20]
port 56 nsew signal output
rlabel metal2 s 61696 297072 61752 297872 6 Do[21]
port 57 nsew signal output
rlabel metal2 s 64640 297072 64696 297872 6 Do[22]
port 58 nsew signal output
rlabel metal2 s 67584 297072 67640 297872 6 Do[23]
port 59 nsew signal output
rlabel metal2 s 70436 297072 70492 297872 6 Do[24]
port 60 nsew signal output
rlabel metal2 s 73380 297072 73436 297872 6 Do[25]
port 61 nsew signal output
rlabel metal2 s 76324 297072 76380 297872 6 Do[26]
port 62 nsew signal output
rlabel metal2 s 79268 297072 79324 297872 6 Do[27]
port 63 nsew signal output
rlabel metal2 s 82212 297072 82268 297872 6 Do[28]
port 64 nsew signal output
rlabel metal2 s 85064 297072 85120 297872 6 Do[29]
port 65 nsew signal output
rlabel metal2 s 6128 297072 6184 297872 6 Do[2]
port 66 nsew signal output
rlabel metal2 s 88008 297072 88064 297872 6 Do[30]
port 67 nsew signal output
rlabel metal2 s 90952 297072 91008 297872 6 Do[31]
port 68 nsew signal output
rlabel metal2 s 9072 297072 9128 297872 6 Do[3]
port 69 nsew signal output
rlabel metal2 s 12016 297072 12072 297872 6 Do[4]
port 70 nsew signal output
rlabel metal2 s 14868 297072 14924 297872 6 Do[5]
port 71 nsew signal output
rlabel metal2 s 17812 297072 17868 297872 6 Do[6]
port 72 nsew signal output
rlabel metal2 s 20756 297072 20812 297872 6 Do[7]
port 73 nsew signal output
rlabel metal2 s 23700 297072 23756 297872 6 Do[8]
port 74 nsew signal output
rlabel metal2 s 26644 297072 26700 297872 6 Do[9]
port 75 nsew signal output
rlabel metal2 s 137780 297072 137836 297872 6 EN
port 76 nsew signal input
rlabel metal2 s 126004 297072 126060 297872 6 WE[0]
port 77 nsew signal input
rlabel metal2 s 128948 297072 129004 297872 6 WE[1]
port 78 nsew signal input
rlabel metal2 s 131892 297072 131948 297872 6 WE[2]
port 79 nsew signal input
rlabel metal2 s 134836 297072 134892 297872 6 WE[3]
port 80 nsew signal input
rlabel metal4 s 219142 0 219462 295488 6 VPWR
port 81 nsew power bidirectional
rlabel metal4 s 195142 0 195462 295488 6 VPWR
port 82 nsew power bidirectional
rlabel metal4 s 171142 0 171462 295488 6 VPWR
port 83 nsew power bidirectional
rlabel metal4 s 147142 0 147462 295488 6 VPWR
port 84 nsew power bidirectional
rlabel metal4 s 123142 0 123462 295488 6 VPWR
port 85 nsew power bidirectional
rlabel metal4 s 99142 0 99462 295488 6 VPWR
port 86 nsew power bidirectional
rlabel metal4 s 75142 0 75462 295488 6 VPWR
port 87 nsew power bidirectional
rlabel metal4 s 51142 0 51462 295488 6 VPWR
port 88 nsew power bidirectional
rlabel metal4 s 27142 0 27462 295488 6 VPWR
port 89 nsew power bidirectional
rlabel metal4 s 3142 0 3462 295488 6 VPWR
port 90 nsew power bidirectional
rlabel metal4 s 231142 0 231462 295488 6 VGND
port 91 nsew ground bidirectional
rlabel metal4 s 207142 0 207462 295488 6 VGND
port 92 nsew ground bidirectional
rlabel metal4 s 183142 0 183462 295488 6 VGND
port 93 nsew ground bidirectional
rlabel metal4 s 159142 0 159462 295488 6 VGND
port 94 nsew ground bidirectional
rlabel metal4 s 135142 0 135462 295488 6 VGND
port 95 nsew ground bidirectional
rlabel metal4 s 111142 0 111462 295488 6 VGND
port 96 nsew ground bidirectional
rlabel metal4 s 87142 0 87462 295488 6 VGND
port 97 nsew ground bidirectional
rlabel metal4 s 63142 0 63462 295488 6 VGND
port 98 nsew ground bidirectional
rlabel metal4 s 39142 0 39462 295488 6 VGND
port 99 nsew ground bidirectional
rlabel metal4 s 15142 0 15462 295488 6 VGND
port 100 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 231824 297872
string LEFview TRUE
<< end >>
