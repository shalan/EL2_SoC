magic
tech sky130A
magscale 1 2
timestamp 1611160305
<< obsli1 >>
rect 1104 1369 138983 77529
<< obsm1 >>
rect 1104 612 138995 78388
<< metal2 >>
rect 70030 78920 70086 79720
<< obsm2 >>
rect 1398 78864 69974 79657
rect 70142 78864 138442 79657
rect 1398 159 138442 78864
<< metal3 >>
rect 139200 79288 140000 79408
rect 139200 78608 140000 78728
rect 0 78064 800 78184
rect 139200 77928 140000 78048
rect 139200 77248 140000 77368
rect 139200 76568 140000 76688
rect 139200 75888 140000 76008
rect 139200 75208 140000 75328
rect 0 74936 800 75056
rect 139200 74528 140000 74648
rect 139200 73848 140000 73968
rect 139200 73168 140000 73288
rect 139200 72488 140000 72608
rect 0 71944 800 72064
rect 139200 71808 140000 71928
rect 139200 71128 140000 71248
rect 139200 70448 140000 70568
rect 139200 69768 140000 69888
rect 139200 69088 140000 69208
rect 0 68816 800 68936
rect 139200 68544 140000 68664
rect 139200 67864 140000 67984
rect 139200 67184 140000 67304
rect 139200 66504 140000 66624
rect 0 65688 800 65808
rect 139200 65824 140000 65944
rect 139200 65144 140000 65264
rect 139200 64464 140000 64584
rect 139200 63784 140000 63904
rect 139200 63104 140000 63224
rect 0 62696 800 62816
rect 139200 62424 140000 62544
rect 139200 61744 140000 61864
rect 139200 61064 140000 61184
rect 139200 60384 140000 60504
rect 0 59568 800 59688
rect 139200 59704 140000 59824
rect 139200 59024 140000 59144
rect 139200 58344 140000 58464
rect 139200 57664 140000 57784
rect 139200 57120 140000 57240
rect 0 56576 800 56696
rect 139200 56440 140000 56560
rect 139200 55760 140000 55880
rect 139200 55080 140000 55200
rect 139200 54400 140000 54520
rect 139200 53720 140000 53840
rect 0 53448 800 53568
rect 139200 53040 140000 53160
rect 139200 52360 140000 52480
rect 139200 51680 140000 51800
rect 139200 51000 140000 51120
rect 0 50320 800 50440
rect 139200 50320 140000 50440
rect 139200 49640 140000 49760
rect 139200 48960 140000 49080
rect 139200 48280 140000 48400
rect 139200 47600 140000 47720
rect 0 47328 800 47448
rect 139200 46920 140000 47040
rect 139200 46240 140000 46360
rect 139200 45696 140000 45816
rect 139200 45016 140000 45136
rect 0 44200 800 44320
rect 139200 44336 140000 44456
rect 139200 43656 140000 43776
rect 139200 42976 140000 43096
rect 139200 42296 140000 42416
rect 139200 41616 140000 41736
rect 0 41208 800 41328
rect 139200 40936 140000 41056
rect 139200 40256 140000 40376
rect 139200 39576 140000 39696
rect 139200 38896 140000 39016
rect 0 38080 800 38200
rect 139200 38216 140000 38336
rect 139200 37536 140000 37656
rect 139200 36856 140000 36976
rect 139200 36176 140000 36296
rect 139200 35496 140000 35616
rect 0 34952 800 35072
rect 139200 34816 140000 34936
rect 139200 34272 140000 34392
rect 139200 33592 140000 33712
rect 139200 32912 140000 33032
rect 139200 32232 140000 32352
rect 0 31960 800 32080
rect 139200 31552 140000 31672
rect 139200 30872 140000 30992
rect 139200 30192 140000 30312
rect 139200 29512 140000 29632
rect 0 28832 800 28952
rect 139200 28832 140000 28952
rect 139200 28152 140000 28272
rect 139200 27472 140000 27592
rect 139200 26792 140000 26912
rect 139200 26112 140000 26232
rect 0 25704 800 25824
rect 139200 25432 140000 25552
rect 139200 24752 140000 24872
rect 139200 24072 140000 24192
rect 139200 23392 140000 23512
rect 0 22712 800 22832
rect 139200 22848 140000 22968
rect 139200 22168 140000 22288
rect 139200 21488 140000 21608
rect 139200 20808 140000 20928
rect 139200 20128 140000 20248
rect 0 19584 800 19704
rect 139200 19448 140000 19568
rect 139200 18768 140000 18888
rect 139200 18088 140000 18208
rect 139200 17408 140000 17528
rect 0 16592 800 16712
rect 139200 16728 140000 16848
rect 139200 16048 140000 16168
rect 139200 15368 140000 15488
rect 139200 14688 140000 14808
rect 139200 14008 140000 14128
rect 0 13464 800 13584
rect 139200 13328 140000 13448
rect 139200 12648 140000 12768
rect 139200 11968 140000 12088
rect 139200 11424 140000 11544
rect 139200 10744 140000 10864
rect 0 10336 800 10456
rect 139200 10064 140000 10184
rect 139200 9384 140000 9504
rect 139200 8704 140000 8824
rect 139200 8024 140000 8144
rect 0 7344 800 7464
rect 139200 7344 140000 7464
rect 139200 6664 140000 6784
rect 139200 5984 140000 6104
rect 139200 5304 140000 5424
rect 139200 4624 140000 4744
rect 0 4216 800 4336
rect 139200 3944 140000 4064
rect 139200 3264 140000 3384
rect 139200 2584 140000 2704
rect 139200 1904 140000 2024
rect 0 1224 800 1344
rect 139200 1224 140000 1344
rect 139200 544 140000 664
rect 139200 0 140000 120
<< obsm3 >>
rect 798 79488 139226 79653
rect 798 79208 139120 79488
rect 798 78808 139226 79208
rect 798 78528 139120 78808
rect 798 78264 139226 78528
rect 880 78128 139226 78264
rect 880 77984 139120 78128
rect 798 77848 139120 77984
rect 798 77448 139226 77848
rect 798 77168 139120 77448
rect 798 76768 139226 77168
rect 798 76488 139120 76768
rect 798 76088 139226 76488
rect 798 75808 139120 76088
rect 798 75408 139226 75808
rect 798 75136 139120 75408
rect 880 75128 139120 75136
rect 880 74856 139226 75128
rect 798 74728 139226 74856
rect 798 74448 139120 74728
rect 798 74048 139226 74448
rect 798 73768 139120 74048
rect 798 73368 139226 73768
rect 798 73088 139120 73368
rect 798 72688 139226 73088
rect 798 72408 139120 72688
rect 798 72144 139226 72408
rect 880 72008 139226 72144
rect 880 71864 139120 72008
rect 798 71728 139120 71864
rect 798 71328 139226 71728
rect 798 71048 139120 71328
rect 798 70648 139226 71048
rect 798 70368 139120 70648
rect 798 69968 139226 70368
rect 798 69688 139120 69968
rect 798 69288 139226 69688
rect 798 69016 139120 69288
rect 880 69008 139120 69016
rect 880 68744 139226 69008
rect 880 68736 139120 68744
rect 798 68464 139120 68736
rect 798 68064 139226 68464
rect 798 67784 139120 68064
rect 798 67384 139226 67784
rect 798 67104 139120 67384
rect 798 66704 139226 67104
rect 798 66424 139120 66704
rect 798 66024 139226 66424
rect 798 65888 139120 66024
rect 880 65744 139120 65888
rect 880 65608 139226 65744
rect 798 65344 139226 65608
rect 798 65064 139120 65344
rect 798 64664 139226 65064
rect 798 64384 139120 64664
rect 798 63984 139226 64384
rect 798 63704 139120 63984
rect 798 63304 139226 63704
rect 798 63024 139120 63304
rect 798 62896 139226 63024
rect 880 62624 139226 62896
rect 880 62616 139120 62624
rect 798 62344 139120 62616
rect 798 61944 139226 62344
rect 798 61664 139120 61944
rect 798 61264 139226 61664
rect 798 60984 139120 61264
rect 798 60584 139226 60984
rect 798 60304 139120 60584
rect 798 59904 139226 60304
rect 798 59768 139120 59904
rect 880 59624 139120 59768
rect 880 59488 139226 59624
rect 798 59224 139226 59488
rect 798 58944 139120 59224
rect 798 58544 139226 58944
rect 798 58264 139120 58544
rect 798 57864 139226 58264
rect 798 57584 139120 57864
rect 798 57320 139226 57584
rect 798 57040 139120 57320
rect 798 56776 139226 57040
rect 880 56640 139226 56776
rect 880 56496 139120 56640
rect 798 56360 139120 56496
rect 798 55960 139226 56360
rect 798 55680 139120 55960
rect 798 55280 139226 55680
rect 798 55000 139120 55280
rect 798 54600 139226 55000
rect 798 54320 139120 54600
rect 798 53920 139226 54320
rect 798 53648 139120 53920
rect 880 53640 139120 53648
rect 880 53368 139226 53640
rect 798 53240 139226 53368
rect 798 52960 139120 53240
rect 798 52560 139226 52960
rect 798 52280 139120 52560
rect 798 51880 139226 52280
rect 798 51600 139120 51880
rect 798 51200 139226 51600
rect 798 50920 139120 51200
rect 798 50520 139226 50920
rect 880 50240 139120 50520
rect 798 49840 139226 50240
rect 798 49560 139120 49840
rect 798 49160 139226 49560
rect 798 48880 139120 49160
rect 798 48480 139226 48880
rect 798 48200 139120 48480
rect 798 47800 139226 48200
rect 798 47528 139120 47800
rect 880 47520 139120 47528
rect 880 47248 139226 47520
rect 798 47120 139226 47248
rect 798 46840 139120 47120
rect 798 46440 139226 46840
rect 798 46160 139120 46440
rect 798 45896 139226 46160
rect 798 45616 139120 45896
rect 798 45216 139226 45616
rect 798 44936 139120 45216
rect 798 44536 139226 44936
rect 798 44400 139120 44536
rect 880 44256 139120 44400
rect 880 44120 139226 44256
rect 798 43856 139226 44120
rect 798 43576 139120 43856
rect 798 43176 139226 43576
rect 798 42896 139120 43176
rect 798 42496 139226 42896
rect 798 42216 139120 42496
rect 798 41816 139226 42216
rect 798 41536 139120 41816
rect 798 41408 139226 41536
rect 880 41136 139226 41408
rect 880 41128 139120 41136
rect 798 40856 139120 41128
rect 798 40456 139226 40856
rect 798 40176 139120 40456
rect 798 39776 139226 40176
rect 798 39496 139120 39776
rect 798 39096 139226 39496
rect 798 38816 139120 39096
rect 798 38416 139226 38816
rect 798 38280 139120 38416
rect 880 38136 139120 38280
rect 880 38000 139226 38136
rect 798 37736 139226 38000
rect 798 37456 139120 37736
rect 798 37056 139226 37456
rect 798 36776 139120 37056
rect 798 36376 139226 36776
rect 798 36096 139120 36376
rect 798 35696 139226 36096
rect 798 35416 139120 35696
rect 798 35152 139226 35416
rect 880 35016 139226 35152
rect 880 34872 139120 35016
rect 798 34736 139120 34872
rect 798 34472 139226 34736
rect 798 34192 139120 34472
rect 798 33792 139226 34192
rect 798 33512 139120 33792
rect 798 33112 139226 33512
rect 798 32832 139120 33112
rect 798 32432 139226 32832
rect 798 32160 139120 32432
rect 880 32152 139120 32160
rect 880 31880 139226 32152
rect 798 31752 139226 31880
rect 798 31472 139120 31752
rect 798 31072 139226 31472
rect 798 30792 139120 31072
rect 798 30392 139226 30792
rect 798 30112 139120 30392
rect 798 29712 139226 30112
rect 798 29432 139120 29712
rect 798 29032 139226 29432
rect 880 28752 139120 29032
rect 798 28352 139226 28752
rect 798 28072 139120 28352
rect 798 27672 139226 28072
rect 798 27392 139120 27672
rect 798 26992 139226 27392
rect 798 26712 139120 26992
rect 798 26312 139226 26712
rect 798 26032 139120 26312
rect 798 25904 139226 26032
rect 880 25632 139226 25904
rect 880 25624 139120 25632
rect 798 25352 139120 25624
rect 798 24952 139226 25352
rect 798 24672 139120 24952
rect 798 24272 139226 24672
rect 798 23992 139120 24272
rect 798 23592 139226 23992
rect 798 23312 139120 23592
rect 798 23048 139226 23312
rect 798 22912 139120 23048
rect 880 22768 139120 22912
rect 880 22632 139226 22768
rect 798 22368 139226 22632
rect 798 22088 139120 22368
rect 798 21688 139226 22088
rect 798 21408 139120 21688
rect 798 21008 139226 21408
rect 798 20728 139120 21008
rect 798 20328 139226 20728
rect 798 20048 139120 20328
rect 798 19784 139226 20048
rect 880 19648 139226 19784
rect 880 19504 139120 19648
rect 798 19368 139120 19504
rect 798 18968 139226 19368
rect 798 18688 139120 18968
rect 798 18288 139226 18688
rect 798 18008 139120 18288
rect 798 17608 139226 18008
rect 798 17328 139120 17608
rect 798 16928 139226 17328
rect 798 16792 139120 16928
rect 880 16648 139120 16792
rect 880 16512 139226 16648
rect 798 16248 139226 16512
rect 798 15968 139120 16248
rect 798 15568 139226 15968
rect 798 15288 139120 15568
rect 798 14888 139226 15288
rect 798 14608 139120 14888
rect 798 14208 139226 14608
rect 798 13928 139120 14208
rect 798 13664 139226 13928
rect 880 13528 139226 13664
rect 880 13384 139120 13528
rect 798 13248 139120 13384
rect 798 12848 139226 13248
rect 798 12568 139120 12848
rect 798 12168 139226 12568
rect 798 11888 139120 12168
rect 798 11624 139226 11888
rect 798 11344 139120 11624
rect 798 10944 139226 11344
rect 798 10664 139120 10944
rect 798 10536 139226 10664
rect 880 10264 139226 10536
rect 880 10256 139120 10264
rect 798 9984 139120 10256
rect 798 9584 139226 9984
rect 798 9304 139120 9584
rect 798 8904 139226 9304
rect 798 8624 139120 8904
rect 798 8224 139226 8624
rect 798 7944 139120 8224
rect 798 7544 139226 7944
rect 880 7264 139120 7544
rect 798 6864 139226 7264
rect 798 6584 139120 6864
rect 798 6184 139226 6584
rect 798 5904 139120 6184
rect 798 5504 139226 5904
rect 798 5224 139120 5504
rect 798 4824 139226 5224
rect 798 4544 139120 4824
rect 798 4416 139226 4544
rect 880 4144 139226 4416
rect 880 4136 139120 4144
rect 798 3864 139120 4136
rect 798 3464 139226 3864
rect 798 3184 139120 3464
rect 798 2784 139226 3184
rect 798 2504 139120 2784
rect 798 2104 139226 2504
rect 798 1824 139120 2104
rect 798 1424 139226 1824
rect 880 1144 139120 1424
rect 798 744 139226 1144
rect 798 464 139120 744
rect 798 200 139226 464
rect 798 163 139120 200
<< metal4 >>
rect 4208 1848 4528 77560
rect 19568 1848 19888 77560
rect 34928 1848 35248 77560
rect 50288 1848 50608 77560
rect 65648 1848 65968 77560
rect 81008 1848 81328 77560
rect 96368 1848 96688 77560
rect 111728 1848 112048 77560
rect 127088 1848 127408 77560
<< obsm4 >>
rect 28947 77640 137389 79653
rect 28947 1768 34848 77640
rect 35328 1768 50208 77640
rect 50688 1768 65568 77640
rect 66048 1768 80928 77640
rect 81408 1768 96288 77640
rect 96768 1768 111648 77640
rect 112128 1768 127008 77640
rect 127488 1768 137389 77640
rect 28947 163 137389 1768
<< labels >>
rlabel metal3 s 139200 0 140000 120 6 HADDR[0]
port 1 nsew signal input
rlabel metal3 s 139200 6664 140000 6784 6 HADDR[10]
port 2 nsew signal input
rlabel metal3 s 139200 7344 140000 7464 6 HADDR[11]
port 3 nsew signal input
rlabel metal3 s 139200 8024 140000 8144 6 HADDR[12]
port 4 nsew signal input
rlabel metal3 s 139200 8704 140000 8824 6 HADDR[13]
port 5 nsew signal input
rlabel metal3 s 139200 9384 140000 9504 6 HADDR[14]
port 6 nsew signal input
rlabel metal3 s 139200 10064 140000 10184 6 HADDR[15]
port 7 nsew signal input
rlabel metal3 s 139200 10744 140000 10864 6 HADDR[16]
port 8 nsew signal input
rlabel metal3 s 139200 11424 140000 11544 6 HADDR[17]
port 9 nsew signal input
rlabel metal3 s 139200 11968 140000 12088 6 HADDR[18]
port 10 nsew signal input
rlabel metal3 s 139200 12648 140000 12768 6 HADDR[19]
port 11 nsew signal input
rlabel metal3 s 139200 544 140000 664 6 HADDR[1]
port 12 nsew signal input
rlabel metal3 s 139200 13328 140000 13448 6 HADDR[20]
port 13 nsew signal input
rlabel metal3 s 139200 14008 140000 14128 6 HADDR[21]
port 14 nsew signal input
rlabel metal3 s 139200 14688 140000 14808 6 HADDR[22]
port 15 nsew signal input
rlabel metal3 s 139200 15368 140000 15488 6 HADDR[23]
port 16 nsew signal input
rlabel metal3 s 139200 16048 140000 16168 6 HADDR[24]
port 17 nsew signal input
rlabel metal3 s 139200 16728 140000 16848 6 HADDR[25]
port 18 nsew signal input
rlabel metal3 s 139200 17408 140000 17528 6 HADDR[26]
port 19 nsew signal input
rlabel metal3 s 139200 18088 140000 18208 6 HADDR[27]
port 20 nsew signal input
rlabel metal3 s 139200 18768 140000 18888 6 HADDR[28]
port 21 nsew signal input
rlabel metal3 s 139200 19448 140000 19568 6 HADDR[29]
port 22 nsew signal input
rlabel metal3 s 139200 1224 140000 1344 6 HADDR[2]
port 23 nsew signal input
rlabel metal3 s 139200 20128 140000 20248 6 HADDR[30]
port 24 nsew signal input
rlabel metal3 s 139200 20808 140000 20928 6 HADDR[31]
port 25 nsew signal input
rlabel metal3 s 139200 1904 140000 2024 6 HADDR[3]
port 26 nsew signal input
rlabel metal3 s 139200 2584 140000 2704 6 HADDR[4]
port 27 nsew signal input
rlabel metal3 s 139200 3264 140000 3384 6 HADDR[5]
port 28 nsew signal input
rlabel metal3 s 139200 3944 140000 4064 6 HADDR[6]
port 29 nsew signal input
rlabel metal3 s 139200 4624 140000 4744 6 HADDR[7]
port 30 nsew signal input
rlabel metal3 s 139200 5304 140000 5424 6 HADDR[8]
port 31 nsew signal input
rlabel metal3 s 139200 5984 140000 6104 6 HADDR[9]
port 32 nsew signal input
rlabel metal3 s 139200 67864 140000 67984 6 HCLK
port 33 nsew signal input
rlabel metal3 s 139200 21488 140000 21608 6 HRDATA[0]
port 34 nsew signal output
rlabel metal3 s 139200 28152 140000 28272 6 HRDATA[10]
port 35 nsew signal output
rlabel metal3 s 139200 28832 140000 28952 6 HRDATA[11]
port 36 nsew signal output
rlabel metal3 s 139200 29512 140000 29632 6 HRDATA[12]
port 37 nsew signal output
rlabel metal3 s 139200 30192 140000 30312 6 HRDATA[13]
port 38 nsew signal output
rlabel metal3 s 139200 30872 140000 30992 6 HRDATA[14]
port 39 nsew signal output
rlabel metal3 s 139200 31552 140000 31672 6 HRDATA[15]
port 40 nsew signal output
rlabel metal3 s 139200 32232 140000 32352 6 HRDATA[16]
port 41 nsew signal output
rlabel metal3 s 139200 32912 140000 33032 6 HRDATA[17]
port 42 nsew signal output
rlabel metal3 s 139200 33592 140000 33712 6 HRDATA[18]
port 43 nsew signal output
rlabel metal3 s 139200 34272 140000 34392 6 HRDATA[19]
port 44 nsew signal output
rlabel metal3 s 139200 22168 140000 22288 6 HRDATA[1]
port 45 nsew signal output
rlabel metal3 s 139200 34816 140000 34936 6 HRDATA[20]
port 46 nsew signal output
rlabel metal3 s 139200 35496 140000 35616 6 HRDATA[21]
port 47 nsew signal output
rlabel metal3 s 139200 36176 140000 36296 6 HRDATA[22]
port 48 nsew signal output
rlabel metal3 s 139200 36856 140000 36976 6 HRDATA[23]
port 49 nsew signal output
rlabel metal3 s 139200 37536 140000 37656 6 HRDATA[24]
port 50 nsew signal output
rlabel metal3 s 139200 38216 140000 38336 6 HRDATA[25]
port 51 nsew signal output
rlabel metal3 s 139200 38896 140000 39016 6 HRDATA[26]
port 52 nsew signal output
rlabel metal3 s 139200 39576 140000 39696 6 HRDATA[27]
port 53 nsew signal output
rlabel metal3 s 139200 40256 140000 40376 6 HRDATA[28]
port 54 nsew signal output
rlabel metal3 s 139200 40936 140000 41056 6 HRDATA[29]
port 55 nsew signal output
rlabel metal3 s 139200 22848 140000 22968 6 HRDATA[2]
port 56 nsew signal output
rlabel metal3 s 139200 41616 140000 41736 6 HRDATA[30]
port 57 nsew signal output
rlabel metal3 s 139200 42296 140000 42416 6 HRDATA[31]
port 58 nsew signal output
rlabel metal3 s 139200 23392 140000 23512 6 HRDATA[3]
port 59 nsew signal output
rlabel metal3 s 139200 24072 140000 24192 6 HRDATA[4]
port 60 nsew signal output
rlabel metal3 s 139200 24752 140000 24872 6 HRDATA[5]
port 61 nsew signal output
rlabel metal3 s 139200 25432 140000 25552 6 HRDATA[6]
port 62 nsew signal output
rlabel metal3 s 139200 26112 140000 26232 6 HRDATA[7]
port 63 nsew signal output
rlabel metal3 s 139200 26792 140000 26912 6 HRDATA[8]
port 64 nsew signal output
rlabel metal3 s 139200 27472 140000 27592 6 HRDATA[9]
port 65 nsew signal output
rlabel metal3 s 139200 66504 140000 66624 6 HREADY
port 66 nsew signal input
rlabel metal2 s 70030 78920 70086 79720 6 HREADYOUT
port 67 nsew signal output
rlabel metal3 s 139200 68544 140000 68664 6 HRESETn
port 68 nsew signal input
rlabel metal3 s 139200 67184 140000 67304 6 HSEL
port 69 nsew signal input
rlabel metal3 s 139200 64464 140000 64584 6 HTRANS[0]
port 70 nsew signal input
rlabel metal3 s 139200 65144 140000 65264 6 HTRANS[1]
port 71 nsew signal input
rlabel metal3 s 139200 42976 140000 43096 6 HWDATA[0]
port 72 nsew signal input
rlabel metal3 s 139200 49640 140000 49760 6 HWDATA[10]
port 73 nsew signal input
rlabel metal3 s 139200 50320 140000 50440 6 HWDATA[11]
port 74 nsew signal input
rlabel metal3 s 139200 51000 140000 51120 6 HWDATA[12]
port 75 nsew signal input
rlabel metal3 s 139200 51680 140000 51800 6 HWDATA[13]
port 76 nsew signal input
rlabel metal3 s 139200 52360 140000 52480 6 HWDATA[14]
port 77 nsew signal input
rlabel metal3 s 139200 53040 140000 53160 6 HWDATA[15]
port 78 nsew signal input
rlabel metal3 s 139200 53720 140000 53840 6 HWDATA[16]
port 79 nsew signal input
rlabel metal3 s 139200 54400 140000 54520 6 HWDATA[17]
port 80 nsew signal input
rlabel metal3 s 139200 55080 140000 55200 6 HWDATA[18]
port 81 nsew signal input
rlabel metal3 s 139200 55760 140000 55880 6 HWDATA[19]
port 82 nsew signal input
rlabel metal3 s 139200 43656 140000 43776 6 HWDATA[1]
port 83 nsew signal input
rlabel metal3 s 139200 56440 140000 56560 6 HWDATA[20]
port 84 nsew signal input
rlabel metal3 s 139200 57120 140000 57240 6 HWDATA[21]
port 85 nsew signal input
rlabel metal3 s 139200 57664 140000 57784 6 HWDATA[22]
port 86 nsew signal input
rlabel metal3 s 139200 58344 140000 58464 6 HWDATA[23]
port 87 nsew signal input
rlabel metal3 s 139200 59024 140000 59144 6 HWDATA[24]
port 88 nsew signal input
rlabel metal3 s 139200 59704 140000 59824 6 HWDATA[25]
port 89 nsew signal input
rlabel metal3 s 139200 60384 140000 60504 6 HWDATA[26]
port 90 nsew signal input
rlabel metal3 s 139200 61064 140000 61184 6 HWDATA[27]
port 91 nsew signal input
rlabel metal3 s 139200 61744 140000 61864 6 HWDATA[28]
port 92 nsew signal input
rlabel metal3 s 139200 62424 140000 62544 6 HWDATA[29]
port 93 nsew signal input
rlabel metal3 s 139200 44336 140000 44456 6 HWDATA[2]
port 94 nsew signal input
rlabel metal3 s 139200 63104 140000 63224 6 HWDATA[30]
port 95 nsew signal input
rlabel metal3 s 139200 63784 140000 63904 6 HWDATA[31]
port 96 nsew signal input
rlabel metal3 s 139200 45016 140000 45136 6 HWDATA[3]
port 97 nsew signal input
rlabel metal3 s 139200 45696 140000 45816 6 HWDATA[4]
port 98 nsew signal input
rlabel metal3 s 139200 46240 140000 46360 6 HWDATA[5]
port 99 nsew signal input
rlabel metal3 s 139200 46920 140000 47040 6 HWDATA[6]
port 100 nsew signal input
rlabel metal3 s 139200 47600 140000 47720 6 HWDATA[7]
port 101 nsew signal input
rlabel metal3 s 139200 48280 140000 48400 6 HWDATA[8]
port 102 nsew signal input
rlabel metal3 s 139200 48960 140000 49080 6 HWDATA[9]
port 103 nsew signal input
rlabel metal3 s 139200 65824 140000 65944 6 HWRITE
port 104 nsew signal input
rlabel metal3 s 139200 69088 140000 69208 6 IRQ[0]
port 105 nsew signal output
rlabel metal3 s 139200 75888 140000 76008 6 IRQ[10]
port 106 nsew signal output
rlabel metal3 s 139200 76568 140000 76688 6 IRQ[11]
port 107 nsew signal output
rlabel metal3 s 139200 77248 140000 77368 6 IRQ[12]
port 108 nsew signal output
rlabel metal3 s 139200 77928 140000 78048 6 IRQ[13]
port 109 nsew signal output
rlabel metal3 s 139200 78608 140000 78728 6 IRQ[14]
port 110 nsew signal output
rlabel metal3 s 139200 79288 140000 79408 6 IRQ[15]
port 111 nsew signal output
rlabel metal3 s 139200 69768 140000 69888 6 IRQ[1]
port 112 nsew signal output
rlabel metal3 s 139200 70448 140000 70568 6 IRQ[2]
port 113 nsew signal output
rlabel metal3 s 139200 71128 140000 71248 6 IRQ[3]
port 114 nsew signal output
rlabel metal3 s 139200 71808 140000 71928 6 IRQ[4]
port 115 nsew signal output
rlabel metal3 s 139200 72488 140000 72608 6 IRQ[5]
port 116 nsew signal output
rlabel metal3 s 139200 73168 140000 73288 6 IRQ[6]
port 117 nsew signal output
rlabel metal3 s 139200 73848 140000 73968 6 IRQ[7]
port 118 nsew signal output
rlabel metal3 s 139200 74528 140000 74648 6 IRQ[8]
port 119 nsew signal output
rlabel metal3 s 139200 75208 140000 75328 6 IRQ[9]
port 120 nsew signal output
rlabel metal3 s 0 13464 800 13584 6 MSI_S2
port 121 nsew signal input
rlabel metal3 s 0 25704 800 25824 6 MSI_S3
port 122 nsew signal input
rlabel metal3 s 0 16592 800 16712 6 MSO_S2
port 123 nsew signal output
rlabel metal3 s 0 28832 800 28952 6 MSO_S3
port 124 nsew signal output
rlabel metal3 s 0 1224 800 1344 6 RsRx_S0
port 125 nsew signal input
rlabel metal3 s 0 7344 800 7464 6 RsRx_S1
port 126 nsew signal input
rlabel metal3 s 0 4216 800 4336 6 RsTx_S0
port 127 nsew signal output
rlabel metal3 s 0 10336 800 10456 6 RsTx_S1
port 128 nsew signal output
rlabel metal3 s 0 22712 800 22832 6 SCLK_S2
port 129 nsew signal output
rlabel metal3 s 0 34952 800 35072 6 SCLK_S3
port 130 nsew signal output
rlabel metal3 s 0 19584 800 19704 6 SSn_S2
port 131 nsew signal output
rlabel metal3 s 0 31960 800 32080 6 SSn_S3
port 132 nsew signal output
rlabel metal3 s 0 74936 800 75056 6 pwm_S6
port 133 nsew signal output
rlabel metal3 s 0 78064 800 78184 6 pwm_S7
port 134 nsew signal output
rlabel metal3 s 0 38080 800 38200 6 scl_i_S4
port 135 nsew signal input
rlabel metal3 s 0 56576 800 56696 6 scl_i_S5
port 136 nsew signal input
rlabel metal3 s 0 41208 800 41328 6 scl_o_S4
port 137 nsew signal output
rlabel metal3 s 0 59568 800 59688 6 scl_o_S5
port 138 nsew signal output
rlabel metal3 s 0 44200 800 44320 6 scl_oen_o_S4
port 139 nsew signal output
rlabel metal3 s 0 62696 800 62816 6 scl_oen_o_S5
port 140 nsew signal output
rlabel metal3 s 0 47328 800 47448 6 sda_i_S4
port 141 nsew signal input
rlabel metal3 s 0 65688 800 65808 6 sda_i_S5
port 142 nsew signal input
rlabel metal3 s 0 50320 800 50440 6 sda_o_S4
port 143 nsew signal output
rlabel metal3 s 0 68816 800 68936 6 sda_o_S5
port 144 nsew signal output
rlabel metal3 s 0 53448 800 53568 6 sda_oen_o_S4
port 145 nsew signal output
rlabel metal3 s 0 71944 800 72064 6 sda_oen_o_S5
port 146 nsew signal output
rlabel metal4 s 127088 1848 127408 77560 6 VPWR
port 147 nsew power bidirectional
rlabel metal4 s 96368 1848 96688 77560 6 VPWR
port 148 nsew power bidirectional
rlabel metal4 s 65648 1848 65968 77560 6 VPWR
port 149 nsew power bidirectional
rlabel metal4 s 34928 1848 35248 77560 6 VPWR
port 150 nsew power bidirectional
rlabel metal4 s 4208 1848 4528 77560 6 VPWR
port 151 nsew power bidirectional
rlabel metal4 s 111728 1848 112048 77560 6 VGND
port 152 nsew ground bidirectional
rlabel metal4 s 81008 1848 81328 77560 6 VGND
port 153 nsew ground bidirectional
rlabel metal4 s 50288 1848 50608 77560 6 VGND
port 154 nsew ground bidirectional
rlabel metal4 s 19568 1848 19888 77560 6 VGND
port 155 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 140000 79720
string LEFview TRUE
<< end >>
