* NGSPICE file created from apb_sys_0.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt apb_sys_0 HADDR[0] HADDR[10] HADDR[11] HADDR[12] HADDR[13] HADDR[14] HADDR[15]
+ HADDR[16] HADDR[17] HADDR[18] HADDR[19] HADDR[1] HADDR[20] HADDR[21] HADDR[22] HADDR[23]
+ HADDR[24] HADDR[25] HADDR[26] HADDR[27] HADDR[28] HADDR[29] HADDR[2] HADDR[30] HADDR[31]
+ HADDR[3] HADDR[4] HADDR[5] HADDR[6] HADDR[7] HADDR[8] HADDR[9] HCLK HRDATA[0] HRDATA[10]
+ HRDATA[11] HRDATA[12] HRDATA[13] HRDATA[14] HRDATA[15] HRDATA[16] HRDATA[17] HRDATA[18]
+ HRDATA[19] HRDATA[1] HRDATA[20] HRDATA[21] HRDATA[22] HRDATA[23] HRDATA[24] HRDATA[25]
+ HRDATA[26] HRDATA[27] HRDATA[28] HRDATA[29] HRDATA[2] HRDATA[30] HRDATA[31] HRDATA[3]
+ HRDATA[4] HRDATA[5] HRDATA[6] HRDATA[7] HRDATA[8] HRDATA[9] HREADY HREADYOUT HRESETn
+ HSEL HTRANS[0] HTRANS[1] HWDATA[0] HWDATA[10] HWDATA[11] HWDATA[12] HWDATA[13] HWDATA[14]
+ HWDATA[15] HWDATA[16] HWDATA[17] HWDATA[18] HWDATA[19] HWDATA[1] HWDATA[20] HWDATA[21]
+ HWDATA[22] HWDATA[23] HWDATA[24] HWDATA[25] HWDATA[26] HWDATA[27] HWDATA[28] HWDATA[29]
+ HWDATA[2] HWDATA[30] HWDATA[31] HWDATA[3] HWDATA[4] HWDATA[5] HWDATA[6] HWDATA[7]
+ HWDATA[8] HWDATA[9] HWRITE IRQ[0] IRQ[10] IRQ[11] IRQ[12] IRQ[13] IRQ[14] IRQ[15]
+ IRQ[1] IRQ[2] IRQ[3] IRQ[4] IRQ[5] IRQ[6] IRQ[7] IRQ[8] IRQ[9] MSI_S2 MSI_S3 MSO_S2
+ MSO_S3 RsRx_S0 RsRx_S1 RsTx_S0 RsTx_S1 SCLK_S2 SCLK_S3 SSn_S2 SSn_S3 pwm_S6 pwm_S7
+ scl_i_S4 scl_i_S5 scl_o_S4 scl_o_S5 scl_oen_o_S4 scl_oen_o_S5 sda_i_S4 sda_i_S5
+ sda_o_S4 sda_o_S5 sda_oen_o_S4 sda_oen_o_S5 VPWR VGND
XFILLER_45_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18869_ _18868_/Y _18866_/X _18802_/X _18866_/X VGND VGND VPWR VPWR _23536_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20900_ _20900_/A VGND VGND VPWR VPWR _22587_/B sky130_fd_sc_hd__buf_2
XANTENNA__13615__A _13614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21880_ _15271_/A _21863_/Y _21870_/Y _21879_/X VGND VGND VPWR VPWR _22004_/A sky130_fd_sc_hd__a211o_4
XFILLER_94_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20831_ _20823_/X _20830_/X _13009_/Y _20823_/X VGND VGND VPWR VPWR _20831_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21832__A _20979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22878__B1 _20821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24992__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22342__A2 _20927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20762_ _16817_/A _14015_/A _20736_/A _15642_/X VGND VGND VPWR VPWR _20762_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24921__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23550_ _23493_/CLK _23550_/D VGND VGND VPWR VPWR _23550_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_74_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16557__B1 _16556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13053__C _13053_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18010__A3 _18000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21550__B1 _24812_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22501_ _22501_/A VGND VGND VPWR VPWR _22580_/B sky130_fd_sc_hd__buf_2
XFILLER_39_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24239__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23481_ _25061_/CLK _23481_/D VGND VGND VPWR VPWR _19024_/A sky130_fd_sc_hd__dfxtp_4
X_20693_ _12013_/A _20693_/B VGND VGND VPWR VPWR _20693_/Y sky130_fd_sc_hd__nor2_4
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_5_13_0_HCLK_A clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22432_ _24409_/Q _20821_/X _21642_/X _22431_/X VGND VGND VPWR VPWR _22432_/X sky130_fd_sc_hd__a211o_4
XFILLER_104_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25220_ _25217_/CLK _25220_/D HRESETn VGND VGND VPWR VPWR _11496_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16309__B1 _15828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22363_ _22438_/A _22362_/X VGND VGND VPWR VPWR _22363_/X sky130_fd_sc_hd__and2_4
XANTENNA__12594__B2 _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25151_ _24824_/CLK _11976_/X HRESETn VGND VGND VPWR VPWR _11975_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22382__B _22238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21314_ _24916_/Q _21448_/B VGND VGND VPWR VPWR _21314_/X sky130_fd_sc_hd__and2_4
X_24102_ _24140_/CLK _16662_/X HRESETn VGND VGND VPWR VPWR _14744_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15532__A1 _15430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21279__A _23023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25082_ _25091_/CLK _25082_/D HRESETn VGND VGND VPWR VPWR _25082_/Q sky130_fd_sc_hd__dfrtp_4
X_22294_ _22294_/A _22238_/X VGND VGND VPWR VPWR _22294_/X sky130_fd_sc_hd__or2_4
X_24033_ _24596_/CLK _24033_/D HRESETn VGND VGND VPWR VPWR _16961_/A sky130_fd_sc_hd__dfrtp_4
X_21245_ _22564_/B VGND VGND VPWR VPWR _21245_/X sky130_fd_sc_hd__buf_2
XFILLER_102_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23874__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25098__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21176_ _21149_/X _21174_/X _21175_/X VGND VGND VPWR VPWR _21176_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__20911__A _21357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23803__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25027__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20127_ _20127_/A VGND VGND VPWR VPWR _20127_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20058_ _21649_/C VGND VGND VPWR VPWR _20058_/Y sky130_fd_sc_hd__inv_2
X_24935_ _24974_/CLK _24935_/D HRESETn VGND VGND VPWR VPWR _24935_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11900_ _11900_/A VGND VGND VPWR VPWR _11900_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12880_ _12880_/A _12880_/B _12880_/C _12854_/Y VGND VGND VPWR VPWR _12882_/C sky130_fd_sc_hd__or4_4
XFILLER_2_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24866_ _24870_/CLK _24866_/D HRESETn VGND VGND VPWR VPWR _14059_/A sky130_fd_sc_hd__dfstp_4
XFILLER_22_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_128_0_HCLK clkbuf_7_64_0_HCLK/X VGND VGND VPWR VPWR _24733_/CLK sky130_fd_sc_hd__clkbuf_1
X_11831_ _11830_/Y VGND VGND VPWR VPWR _11831_/X sky130_fd_sc_hd__buf_2
X_23817_ _23824_/CLK _23817_/D HRESETn VGND VGND VPWR VPWR _18419_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_73_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24797_ _24859_/CLK _24797_/D HRESETn VGND VGND VPWR VPWR _14272_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14271__B2 _14268_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14550_ _14548_/X _14549_/X _14548_/X _14549_/X VGND VGND VPWR VPWR _14550_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_54_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24662__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11761_/A _11761_/B _11760_/Y _11761_/Y VGND VGND VPWR VPWR _11763_/D sky130_fd_sc_hd__a211o_4
XFILLER_109_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18001__A3 _18000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23748_ _24180_/CLK _23748_/D HRESETn VGND VGND VPWR VPWR _23748_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13500_/X VGND VGND VPWR VPWR _13501_/Y sky130_fd_sc_hd__inv_2
XPHY_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _21534_/A _14475_/X _14480_/X VGND VGND VPWR VPWR _24752_/D sky130_fd_sc_hd__a21oi_4
X_11693_ _11693_/A _11693_/B _11689_/X _11692_/X VGND VGND VPWR VPWR _11694_/D sky130_fd_sc_hd__or4_4
XPHY_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23679_ _24723_/CLK _20399_/Y HRESETn VGND VGND VPWR VPWR _17183_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _16218_/Y _16138_/A _16219_/X _16138_/A VGND VGND VPWR VPWR _24289_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _13432_/A VGND VGND VPWR VPWR _13432_/Y sky130_fd_sc_hd__inv_2
XPHY_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16151_ _24315_/Q VGND VGND VPWR VPWR _16151_/Y sky130_fd_sc_hd__inv_2
X_13363_ _13363_/A VGND VGND VPWR VPWR _13363_/X sky130_fd_sc_hd__buf_2
X_15102_ _15132_/A _15129_/A VGND VGND VPWR VPWR _15125_/A sky130_fd_sc_hd__or2_4
X_12314_ _12412_/D VGND VGND VPWR VPWR _12474_/C sky130_fd_sc_hd__buf_2
X_16082_ _24340_/Q VGND VGND VPWR VPWR _16082_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13294_ _13166_/A _20007_/A VGND VGND VPWR VPWR _13295_/C sky130_fd_sc_hd__or2_4
XFILLER_138_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15033_ _15033_/A _15020_/X VGND VGND VPWR VPWR _15034_/B sky130_fd_sc_hd__or2_4
X_19910_ _19910_/A VGND VGND VPWR VPWR _21787_/B sky130_fd_sc_hd__inv_2
X_12245_ _12227_/X _12245_/B _12245_/C VGND VGND VPWR VPWR _25120_/D sky130_fd_sc_hd__and3_4
XFILLER_5_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12176_ _12176_/A _12097_/Y _12103_/Y _12157_/Y VGND VGND VPWR VPWR _12176_/X sky130_fd_sc_hd__or4_4
X_19841_ _19841_/A VGND VGND VPWR VPWR _19841_/X sky130_fd_sc_hd__buf_2
XANTENNA__15287__B1 _15286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20821__A _22148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15915__A _16228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16984_ _24056_/Q VGND VGND VPWR VPWR _17022_/A sky130_fd_sc_hd__inv_2
X_19772_ _19759_/Y VGND VGND VPWR VPWR _19772_/X sky130_fd_sc_hd__buf_2
XFILLER_111_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22021__A1 _22011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15935_ _22838_/A VGND VGND VPWR VPWR _15935_/Y sky130_fd_sc_hd__inv_2
X_18723_ _23586_/Q VGND VGND VPWR VPWR _18723_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_24_0_HCLK clkbuf_6_12_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_24_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19973__B1 _19445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18654_ _18654_/A VGND VGND VPWR VPWR _21508_/B sky130_fd_sc_hd__inv_2
X_15866_ _24411_/Q VGND VGND VPWR VPWR _15866_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_87_0_HCLK clkbuf_7_87_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_87_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14817_ _24690_/Q _24133_/Q _15067_/B _14816_/Y VGND VGND VPWR VPWR _14817_/X sky130_fd_sc_hd__o22a_4
X_17605_ _17603_/A _17605_/B _17605_/C VGND VGND VPWR VPWR _23949_/D sky130_fd_sc_hd__and3_4
X_18585_ _16378_/A _18427_/A _16371_/A _18543_/A VGND VGND VPWR VPWR _18585_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15797_ _15797_/A VGND VGND VPWR VPWR _15797_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17536_ _17482_/A _17535_/Y VGND VGND VPWR VPWR _17538_/B sky130_fd_sc_hd__or2_4
XANTENNA__15650__A _11944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14748_ _24684_/Q _14747_/A _15087_/A _14747_/Y VGND VGND VPWR VPWR _14748_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12273__B1 _12195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17200__B2 _17198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24332__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17467_ _21805_/A _17453_/X _17466_/A _17452_/A VGND VGND VPWR VPWR _17468_/A sky130_fd_sc_hd__o22a_4
X_14679_ _14622_/X _14678_/Y _24867_/Q _14622_/X VGND VGND VPWR VPWR _24718_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14266__A _13934_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16418_ _24212_/Q VGND VGND VPWR VPWR _16418_/Y sky130_fd_sc_hd__inv_2
X_19206_ _19206_/A VGND VGND VPWR VPWR _19206_/Y sky130_fd_sc_hd__inv_2
X_17398_ _17300_/X VGND VGND VPWR VPWR _17423_/A sky130_fd_sc_hd__buf_2
XANTENNA__22483__A _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19137_ _19137_/A VGND VGND VPWR VPWR _19137_/X sky130_fd_sc_hd__buf_2
XFILLER_118_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16349_ _24237_/Q VGND VGND VPWR VPWR _16349_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16481__A _16493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19068_ _17848_/B VGND VGND VPWR VPWR _19068_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23037__B1 _17224_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18019_ _23901_/Q VGND VGND VPWR VPWR _19531_/A sky130_fd_sc_hd__buf_2
X_21030_ _20783_/X VGND VGND VPWR VPWR _21030_/X sky130_fd_sc_hd__buf_2
XANTENNA__25191__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25120__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22981_ _12391_/Y _22259_/X _17021_/A _22433_/A VGND VGND VPWR VPWR _22982_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12500__A1 _12495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19964__B1 _19963_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24720_ _24723_/CLK _14672_/X HRESETn VGND VGND VPWR VPWR _14625_/A sky130_fd_sc_hd__dfrtp_4
X_21932_ _21342_/A _21932_/B VGND VGND VPWR VPWR _21932_/X sky130_fd_sc_hd__or2_4
XANTENNA__21562__A _21562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24651_ _24654_/CLK _24651_/D HRESETn VGND VGND VPWR VPWR _24651_/Q sky130_fd_sc_hd__dfrtp_4
X_21863_ _21863_/A VGND VGND VPWR VPWR _21863_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23602_ _23992_/CLK _18680_/X VGND VGND VPWR VPWR _23602_/Q sky130_fd_sc_hd__dfxtp_4
X_20814_ _21565_/A VGND VGND VPWR VPWR _20814_/X sky130_fd_sc_hd__buf_2
X_21794_ _21292_/A VGND VGND VPWR VPWR _21868_/B sky130_fd_sc_hd__buf_2
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24582_ _24017_/CLK _15423_/X HRESETn VGND VGND VPWR VPWR _20550_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_24_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24073__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23533_ _23531_/CLK _18881_/X VGND VGND VPWR VPWR _23533_/Q sky130_fd_sc_hd__dfxtp_4
X_20745_ _20744_/X VGND VGND VPWR VPWR _20745_/X sky130_fd_sc_hd__buf_2
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24002__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20676_ _23756_/Q _23755_/Q _13541_/X VGND VGND VPWR VPWR _20676_/X sky130_fd_sc_hd__or3_4
XFILLER_50_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23464_ _23419_/CLK _23464_/D VGND VGND VPWR VPWR _23464_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25203_ _23969_/CLK _25203_/D HRESETn VGND VGND VPWR VPWR _11587_/A sky130_fd_sc_hd__dfrtp_4
X_22415_ _22414_/X VGND VGND VPWR VPWR _22416_/D sky130_fd_sc_hd__inv_2
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16391__A _21109_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23395_ _23411_/CLK _19269_/X VGND VGND VPWR VPWR _21701_/D sky130_fd_sc_hd__dfxtp_4
X_25134_ _25141_/CLK _25134_/D HRESETn VGND VGND VPWR VPWR _12069_/A sky130_fd_sc_hd__dfrtp_4
X_22346_ _21529_/X _22342_/X _22500_/A _22345_/X VGND VGND VPWR VPWR _22346_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25208__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22277_ _22512_/A VGND VGND VPWR VPWR _22495_/A sky130_fd_sc_hd__buf_2
X_25065_ _25046_/CLK _12676_/Y HRESETn VGND VGND VPWR VPWR _25065_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23043__A3 HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12030_ _23796_/Q _12015_/B _12029_/Y VGND VGND VPWR VPWR _20696_/A sky130_fd_sc_hd__o21a_4
XANTENNA__17258__A1 _25197_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21228_ _21234_/A VGND VGND VPWR VPWR _21229_/A sky130_fd_sc_hd__buf_2
X_24016_ _24017_/CLK _24016_/D HRESETn VGND VGND VPWR VPWR _17208_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15735__A _15431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21159_ _21159_/A _19661_/Y VGND VGND VPWR VPWR _21160_/C sky130_fd_sc_hd__or2_4
XFILLER_8_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13981_ _13981_/A VGND VGND VPWR VPWR _13981_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15720_ _15720_/A VGND VGND VPWR VPWR _15720_/X sky130_fd_sc_hd__buf_2
X_12932_ _12932_/A VGND VGND VPWR VPWR _12932_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17950__A _17918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24918_ _24923_/CLK _13701_/X HRESETn VGND VGND VPWR VPWR _24918_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24843__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15651_ _15421_/X _15647_/X _15635_/X _24499_/Q _15650_/X VGND VGND VPWR VPWR _24499_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_98_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12863_ _25011_/Q VGND VGND VPWR VPWR _12863_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19292__A2_N _19289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24849_ _24840_/CLK _14124_/Y HRESETn VGND VGND VPWR VPWR _11917_/D sky130_fd_sc_hd__dfrtp_4
XANTENNA__16566__A _16566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14602_ _19946_/A _19946_/B VGND VGND VPWR VPWR _19167_/B sky130_fd_sc_hd__or2_4
XANTENNA__15470__A _15464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11814_ _11817_/B VGND VGND VPWR VPWR _11814_/Y sky130_fd_sc_hd__inv_2
X_18370_ _23842_/Q VGND VGND VPWR VPWR _18412_/A sky130_fd_sc_hd__inv_2
X_15582_ _15582_/A VGND VGND VPWR VPWR _15582_/X sky130_fd_sc_hd__buf_2
XANTENNA__22718__D _22718_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12794_ _12793_/Y _20834_/A _12793_/Y _20834_/A VGND VGND VPWR VPWR _12795_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _23982_/Q VGND VGND VPWR VPWR _17321_/Y sky130_fd_sc_hd__inv_2
X_14533_ _20994_/A VGND VGND VPWR VPWR _21009_/A sky130_fd_sc_hd__buf_2
XFILLER_30_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11745_/A _11745_/B VGND VGND VPWR VPWR _11763_/C sky130_fd_sc_hd__or2_4
XFILLER_30_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11503__A _11503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _11565_/A _17251_/A _11565_/Y _17251_/Y VGND VGND VPWR VPWR _17252_/X sky130_fd_sc_hd__o22a_4
X_14464_ _14541_/D VGND VGND VPWR VPWR _19779_/B sky130_fd_sc_hd__inv_2
XPHY_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _11676_/A VGND VGND VPWR VPWR _11676_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ _16196_/A VGND VGND VPWR VPWR _16203_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13415_ _24931_/Q VGND VGND VPWR VPWR _13415_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12558__B2 _24528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17183_ _17183_/A _20394_/A VGND VGND VPWR VPWR _17186_/B sky130_fd_sc_hd__or2_4
X_14395_ _14387_/C _14392_/X VGND VGND VPWR VPWR _14395_/X sky130_fd_sc_hd__or2_4
XANTENNA__23796__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16134_ _15655_/A VGND VGND VPWR VPWR _16134_/X sky130_fd_sc_hd__buf_2
X_13346_ _24991_/Q VGND VGND VPWR VPWR _13346_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23725__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16065_ _16063_/Y _16059_/X _15761_/X _16064_/X VGND VGND VPWR VPWR _24348_/D sky130_fd_sc_hd__a2bb2o_4
X_13277_ _13309_/A _13277_/B VGND VGND VPWR VPWR _13278_/C sky130_fd_sc_hd__or2_4
XANTENNA__12334__A _25077_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15016_ _15016_/A _15013_/B _15015_/X VGND VGND VPWR VPWR _15017_/A sky130_fd_sc_hd__or3_4
XFILLER_64_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12228_ _12167_/Y _12183_/B VGND VGND VPWR VPWR _12228_/X sky130_fd_sc_hd__or2_4
XANTENNA__22793__A2 _20757_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19824_ _23195_/Q VGND VGND VPWR VPWR _19824_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15645__A _15459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12159_ _12157_/Y _12075_/A _12265_/A _24548_/Q VGND VGND VPWR VPWR _12159_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19245__A2_N _19239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19755_ _25169_/Q VGND VGND VPWR VPWR _19755_/X sky130_fd_sc_hd__buf_2
X_16967_ _16193_/A _16966_/Y _16151_/Y _24053_/Q VGND VGND VPWR VPWR _16972_/B sky130_fd_sc_hd__a2bb2o_4
X_18706_ _16291_/A VGND VGND VPWR VPWR _18706_/X sky130_fd_sc_hd__buf_2
X_15918_ _23002_/A VGND VGND VPWR VPWR _15918_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24584__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16898_ _16823_/Y _16898_/B VGND VGND VPWR VPWR _16902_/B sky130_fd_sc_hd__or2_4
X_19686_ _23246_/Q VGND VGND VPWR VPWR _19686_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15849_ _15849_/A VGND VGND VPWR VPWR _15849_/Y sky130_fd_sc_hd__inv_2
X_18637_ _11701_/C VGND VGND VPWR VPWR _18637_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24513__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_111_0_HCLK clkbuf_7_55_0_HCLK/X VGND VGND VPWR VPWR _24349_/CLK sky130_fd_sc_hd__clkbuf_1
X_18568_ _16387_/Y _18355_/X _16387_/Y _18355_/X VGND VGND VPWR VPWR _18568_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_174_0_HCLK clkbuf_7_87_0_HCLK/X VGND VGND VPWR VPWR _23303_/CLK sky130_fd_sc_hd__clkbuf_1
X_17519_ _17509_/A _17517_/X _17519_/C VGND VGND VPWR VPWR _23971_/D sky130_fd_sc_hd__and3_4
X_18499_ _18495_/B _18502_/A VGND VGND VPWR VPWR _18504_/B sky130_fd_sc_hd__or2_4
XFILLER_127_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18691__A _18690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20530_ _20511_/X _20529_/X _15339_/A _20515_/X VGND VGND VPWR VPWR _20530_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14538__A2 _14521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20461_ _20511_/A VGND VGND VPWR VPWR _20461_/X sky130_fd_sc_hd__buf_2
X_22200_ _22191_/X _22194_/Y _22167_/A _22199_/X VGND VGND VPWR VPWR _22200_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23180_ _23154_/CLK _23180_/D VGND VGND VPWR VPWR _19868_/A sky130_fd_sc_hd__dfxtp_4
X_20392_ _20391_/X VGND VGND VPWR VPWR _20392_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22131_ _22129_/X _22130_/X _21994_/X _24552_/Q _21995_/X VGND VGND VPWR VPWR _22131_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_47_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22062_ _21675_/A _22060_/X _22061_/X VGND VGND VPWR VPWR _22066_/B sky130_fd_sc_hd__and3_4
XANTENNA__14783__A2_N _14781_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22233__A1 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22233__B2 _22228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20461__A _20511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21013_ _20994_/A _21013_/B VGND VGND VPWR VPWR _21013_/X sky130_fd_sc_hd__or2_4
XANTENNA__22784__A2 _20821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20795__A1 _25190_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19937__B1 _19455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15671__B1 _24493_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22964_ _22955_/X _22959_/X _22964_/C VGND VGND VPWR VPWR _22964_/X sky130_fd_sc_hd__or3_4
XANTENNA__21292__A _21292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24703_ _24706_/CLK _24703_/D HRESETn VGND VGND VPWR VPWR _14874_/A sky130_fd_sc_hd__dfrtp_4
X_21915_ _21930_/A _21911_/X _21914_/X VGND VGND VPWR VPWR _21915_/X sky130_fd_sc_hd__or3_4
XANTENNA__24254__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_70_0_HCLK clkbuf_7_71_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_70_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22895_ _21572_/B _22894_/X _22640_/X _25217_/Q _22641_/X VGND VGND VPWR VPWR _22895_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15423__B1 _20550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24634_ _24641_/CLK _15268_/X HRESETn VGND VGND VPWR VPWR _13754_/A sky130_fd_sc_hd__dfrtp_4
X_21846_ _21042_/A _21845_/X _21432_/C _24550_/Q _20900_/A VGND VGND VPWR VPWR _21847_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24565_ _24573_/CLK _24565_/D HRESETn VGND VGND VPWR VPWR _24565_/Q sky130_fd_sc_hd__dfrtp_4
X_21777_ _21777_/A _21777_/B VGND VGND VPWR VPWR _21777_/X sky130_fd_sc_hd__or2_4
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11530_ _22992_/B VGND VGND VPWR VPWR _11530_/X sky130_fd_sc_hd__buf_2
XFILLER_11_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23516_ _23514_/CLK _23516_/D VGND VGND VPWR VPWR _18926_/A sky130_fd_sc_hd__dfxtp_4
X_20728_ _20729_/A _23665_/D _23666_/Q VGND VGND VPWR VPWR _20728_/X sky130_fd_sc_hd__and3_4
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24496_ _24604_/CLK _15667_/X HRESETn VGND VGND VPWR VPWR _24496_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23012__A _23012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23447_ _23425_/CLK _19121_/X VGND VGND VPWR VPWR _23447_/Q sky130_fd_sc_hd__dfxtp_4
X_20659_ _20658_/X VGND VGND VPWR VPWR _23750_/D sky130_fd_sc_hd__inv_2
XFILLER_104_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13200_ _13232_/A _13196_/X _13200_/C VGND VGND VPWR VPWR _13200_/X sky130_fd_sc_hd__or3_4
XFILLER_137_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14180_ _14150_/X VGND VGND VPWR VPWR _14180_/X sky130_fd_sc_hd__buf_2
XFILLER_99_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18676__B1 _16546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23378_ _25002_/CLK _19317_/X VGND VGND VPWR VPWR _23378_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25042__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13131_ _13085_/A _23204_/Q VGND VGND VPWR VPWR _13131_/X sky130_fd_sc_hd__or2_4
X_25117_ _25123_/CLK _25117_/D HRESETn VGND VGND VPWR VPWR _25117_/Q sky130_fd_sc_hd__dfrtp_4
X_22329_ _22175_/A _22327_/X _22349_/B _22328_/X VGND VGND VPWR VPWR _22330_/A sky130_fd_sc_hd__o22a_4
XFILLER_124_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13062_ _13078_/A VGND VGND VPWR VPWR _13202_/A sky130_fd_sc_hd__buf_2
XANTENNA__21467__A _21333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25048_ _25067_/CLK _25048_/D HRESETn VGND VGND VPWR VPWR _25048_/Q sky130_fd_sc_hd__dfrtp_4
X_12013_ _12013_/A _23794_/Q VGND VGND VPWR VPWR _12014_/B sky130_fd_sc_hd__and2_4
XANTENNA__15465__A _15464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17870_ _17934_/A _17870_/B VGND VGND VPWR VPWR _17872_/B sky130_fd_sc_hd__or2_4
XFILLER_117_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16821_ _16821_/A VGND VGND VPWR VPWR _16822_/A sky130_fd_sc_hd__inv_2
XFILLER_78_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19928__B1 _19442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16752_ _15818_/Y _16846_/A _15818_/Y _16846_/A VGND VGND VPWR VPWR _16756_/B sky130_fd_sc_hd__a2bb2o_4
X_19540_ _19538_/Y _19534_/X _11844_/X _19539_/X VGND VGND VPWR VPWR _19540_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13964_ _13937_/X _13962_/X _14255_/A _13963_/X VGND VGND VPWR VPWR _13964_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_93_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15703_ _12357_/Y _15702_/X _15393_/X _15702_/X VGND VGND VPWR VPWR _15703_/X sky130_fd_sc_hd__a2bb2o_4
X_12915_ _12845_/Y _12883_/X _12915_/C VGND VGND VPWR VPWR _12916_/B sky130_fd_sc_hd__or3_4
X_16683_ _15972_/Y _22307_/A _15972_/Y _22307_/A VGND VGND VPWR VPWR _16683_/X sky130_fd_sc_hd__a2bb2o_4
X_19471_ _19470_/Y _19468_/X _19421_/X _19468_/X VGND VGND VPWR VPWR _23325_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25136__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13895_ _13866_/B _13892_/X _13884_/X _13828_/D _13893_/X VGND VGND VPWR VPWR _24910_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_111_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15634_ _12595_/Y _15593_/A _14304_/X _15593_/A VGND VGND VPWR VPWR _15634_/X sky130_fd_sc_hd__a2bb2o_4
X_18422_ _23816_/Q VGND VGND VPWR VPWR _18422_/Y sky130_fd_sc_hd__inv_2
X_12846_ _12845_/Y _12853_/A _22258_/A _12787_/Y VGND VGND VPWR VPWR _12856_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18353_ _23840_/Q VGND VGND VPWR VPWR _18413_/A sky130_fd_sc_hd__inv_2
XANTENNA__21930__A _21930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13976__B1 _24801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15565_ _19859_/A VGND VGND VPWR VPWR _15565_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_247_0_HCLK clkbuf_8_247_0_HCLK/A VGND VGND VPWR VPWR _24681_/CLK sky130_fd_sc_hd__clkbuf_1
X_12777_ _12890_/A _24460_/Q _12890_/A _24460_/Q VGND VGND VPWR VPWR _12783_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23977__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17304_ _17303_/Y VGND VGND VPWR VPWR _17329_/A sky130_fd_sc_hd__buf_2
XFILLER_14_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22745__B _22745_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14508_/X _14515_/Y _24749_/Q _14507_/Y VGND VGND VPWR VPWR _14516_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _11507_/X _11720_/X _11728_/C _11960_/A VGND VGND VPWR VPWR _11728_/X sky130_fd_sc_hd__or4_4
X_18284_ _18284_/A _18277_/X _18283_/Y VGND VGND VPWR VPWR _18284_/X sky130_fd_sc_hd__and3_4
X_15496_ _15482_/X _15483_/X _15494_/X _24561_/Q _15495_/X VGND VGND VPWR VPWR _24561_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23906__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17235_ _17234_/X VGND VGND VPWR VPWR _17235_/Y sky130_fd_sc_hd__inv_2
XPHY_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14447_ _14446_/X VGND VGND VPWR VPWR _14448_/B sky130_fd_sc_hd__inv_2
XFILLER_31_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11659_ _13559_/A _21871_/A _13549_/A _22484_/A VGND VGND VPWR VPWR _11659_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17166_ _17160_/A _17160_/B VGND VGND VPWR VPWR _17166_/Y sky130_fd_sc_hd__nand2_4
X_14378_ _14378_/A VGND VGND VPWR VPWR _14378_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18131__A2 _17052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16117_ _16083_/A VGND VGND VPWR VPWR _16117_/X sky130_fd_sc_hd__buf_2
XFILLER_115_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13329_ _15422_/A _13328_/X VGND VGND VPWR VPWR _13329_/Y sky130_fd_sc_hd__nor2_4
X_17097_ _17097_/A _17097_/B VGND VGND VPWR VPWR _17097_/X sky130_fd_sc_hd__or2_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12064__A _12063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16142__B2 _16138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16048_ _16048_/A VGND VGND VPWR VPWR _16048_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15496__A3 _15494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21377__A _21214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24765__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19807_ _19800_/X _18067_/A _18000_/X _13205_/B _19802_/X VGND VGND VPWR VPWR _23202_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_85_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17999_ _17999_/A VGND VGND VPWR VPWR _17999_/X sky130_fd_sc_hd__buf_2
XFILLER_84_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19919__B1 _19832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19738_ _19737_/Y VGND VGND VPWR VPWR _19738_/X sky130_fd_sc_hd__buf_2
XFILLER_49_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21726__B1 _11532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15822__B _15821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19669_ _22085_/B _19668_/X _19597_/X _19668_/X VGND VGND VPWR VPWR _19669_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_6_57_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21700_ _21700_/A _21756_/B VGND VGND VPWR VPWR _21700_/X sky130_fd_sc_hd__and2_4
XFILLER_53_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22680_ _24565_/Q _22557_/X _22558_/X _22679_/X VGND VGND VPWR VPWR _22681_/C sky130_fd_sc_hd__a211o_4
XANTENNA__21840__A _21840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19147__B2 _19146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21631_ _22084_/A _21631_/B VGND VGND VPWR VPWR _21631_/X sky130_fd_sc_hd__or2_4
XANTENNA__16934__A _16936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24350_ _23872_/CLK _16060_/X HRESETn VGND VGND VPWR VPWR _24350_/Q sky130_fd_sc_hd__dfrtp_4
X_21562_ _21562_/A VGND VGND VPWR VPWR _21562_/X sky130_fd_sc_hd__buf_2
XFILLER_100_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23301_ _23100_/CLK _23301_/D VGND VGND VPWR VPWR _23301_/Q sky130_fd_sc_hd__dfxtp_4
X_20513_ _20512_/A _20513_/B _20517_/A _13497_/D VGND VGND VPWR VPWR _20513_/X sky130_fd_sc_hd__or4_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21493_ _22018_/B _21492_/X _23908_/Q _11941_/X VGND VGND VPWR VPWR _21493_/X sky130_fd_sc_hd__o22a_4
X_24281_ _24104_/CLK _16249_/X HRESETn VGND VGND VPWR VPWR _24281_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22025__A2_N _20818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20444_ _21888_/A _20437_/X _20425_/X _20443_/Y VGND VGND VPWR VPWR _20445_/A sky130_fd_sc_hd__o22a_4
XANTENNA__22454__A1 _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23232_ _23401_/CLK _19732_/X VGND VGND VPWR VPWR _19730_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22454__B2 _22453_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20375_ _15290_/Y _20367_/X _20358_/X _20374_/X VGND VGND VPWR VPWR _20375_/X sky130_fd_sc_hd__a211o_4
X_23163_ _23332_/CLK _23163_/D VGND VGND VPWR VPWR _23163_/Q sky130_fd_sc_hd__dfxtp_4
X_22114_ _11532_/A _20940_/X _22114_/C _22113_/X VGND VGND VPWR VPWR _22114_/X sky130_fd_sc_hd__or4_4
XANTENNA__22206__B2 _22879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23094_ _23383_/CLK _20094_/X VGND VGND VPWR VPWR _23094_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_133_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20191__A _13908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24626__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22045_ _21490_/X _22045_/B _22044_/X VGND VGND VPWR VPWR _22045_/X sky130_fd_sc_hd__and3_4
XFILLER_114_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24435__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23996_ _25214_/CLK _17388_/X HRESETn VGND VGND VPWR VPWR _23996_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22947_ _22946_/X VGND VGND VPWR VPWR _22965_/B sky130_fd_sc_hd__inv_2
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21193__A1 _21176_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12700_ _12700_/A _12700_/B VGND VGND VPWR VPWR _12701_/B sky130_fd_sc_hd__or2_4
X_13680_ _20201_/C _13677_/X _13678_/X _13679_/Y VGND VGND VPWR VPWR _24924_/D sky130_fd_sc_hd__a211o_4
XFILLER_71_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11681__B2 _11680_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22878_ _24152_/Q _22505_/X _20821_/X _22877_/X VGND VGND VPWR VPWR _22879_/C sky130_fd_sc_hd__a211o_4
XFILLER_43_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12631_ _12624_/X _12626_/X _12627_/X _12630_/X VGND VGND VPWR VPWR _12631_/X sky130_fd_sc_hd__or4_4
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24617_ _24618_/CLK _24617_/D HRESETn VGND VGND VPWR VPWR _11499_/A sky130_fd_sc_hd__dfrtp_4
X_21829_ _21825_/X _21828_/X _21172_/X VGND VGND VPWR VPWR _21829_/Y sky130_fd_sc_hd__o21ai_4
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22142__B1 _11954_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22565__B _15655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ HWDATA[21] VGND VGND VPWR VPWR _15350_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_0_0_HCLK clkbuf_6_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12562_ _12562_/A VGND VGND VPWR VPWR _12651_/D sky130_fd_sc_hd__inv_2
XANTENNA__22693__A1 _24345_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24548_ _25084_/CLK _15523_/X HRESETn VGND VGND VPWR VPWR _24548_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_14_0_HCLK clkbuf_7_7_0_HCLK/X VGND VGND VPWR VPWR _23356_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14301_ _14299_/Y _14300_/X _14213_/X _14300_/X VGND VGND VPWR VPWR _24786_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11513_ _24620_/Q _16038_/B _11512_/Y VGND VGND VPWR VPWR _14020_/A sky130_fd_sc_hd__or3_4
XANTENNA__11988__A _21564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15281_ _24628_/Q VGND VGND VPWR VPWR _15281_/Y sky130_fd_sc_hd__inv_2
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _12399_/A VGND VGND VPWR VPWR _12509_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_77_0_HCLK clkbuf_8_77_0_HCLK/A VGND VGND VPWR VPWR _24788_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24479_ _24478_/CLK _24479_/D HRESETn VGND VGND VPWR VPWR _22373_/A sky130_fd_sc_hd__dfrtp_4
X_17020_ _17086_/A VGND VGND VPWR VPWR _17052_/A sky130_fd_sc_hd__buf_2
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14232_ _16373_/A VGND VGND VPWR VPWR _14232_/X sky130_fd_sc_hd__buf_2
XFILLER_138_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22581__A _22351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14163_ _14159_/Y _14155_/X VGND VGND VPWR VPWR _14168_/A sky130_fd_sc_hd__or2_4
X_13114_ _11708_/X VGND VGND VPWR VPWR _13114_/X sky130_fd_sc_hd__buf_2
XFILLER_4_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15478__A3 _15477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14094_ _13398_/A VGND VGND VPWR VPWR _14094_/X sky130_fd_sc_hd__buf_2
X_18971_ _18966_/Y _18970_/X _18901_/X _18970_/X VGND VGND VPWR VPWR _18971_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15883__B1 _15788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13045_ _13045_/A _23076_/Q VGND VGND VPWR VPWR _13045_/X sky130_fd_sc_hd__or2_4
X_17922_ _17725_/A _17922_/B _17922_/C VGND VGND VPWR VPWR _17923_/C sky130_fd_sc_hd__or3_4
XANTENNA__19074__B1 _18938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21925__A _21342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21420__A2 _22154_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24176__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17853_ _17853_/A _23426_/Q VGND VGND VPWR VPWR _17853_/X sky130_fd_sc_hd__or2_4
XFILLER_66_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16804_ _16804_/A _16804_/B _16801_/X _16803_/X VGND VGND VPWR VPWR _16804_/X sky130_fd_sc_hd__or4_4
XFILLER_130_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24105__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21644__B _21181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14996_ _14995_/X VGND VGND VPWR VPWR _14997_/B sky130_fd_sc_hd__inv_2
X_17784_ _17738_/A _17784_/B _17783_/X VGND VGND VPWR VPWR _17785_/C sky130_fd_sc_hd__or3_4
X_19523_ _19510_/Y VGND VGND VPWR VPWR _19523_/X sky130_fd_sc_hd__buf_2
XFILLER_47_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13947_ _13947_/A _13946_/X VGND VGND VPWR VPWR _13947_/Y sky130_fd_sc_hd__nor2_4
X_16735_ _23962_/Q VGND VGND VPWR VPWR _17497_/D sky130_fd_sc_hd__inv_2
XFILLER_75_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16666_ _16643_/A VGND VGND VPWR VPWR _16666_/X sky130_fd_sc_hd__buf_2
X_19454_ _23330_/Q VGND VGND VPWR VPWR _21501_/B sky130_fd_sc_hd__inv_2
X_13878_ _13854_/X _14357_/C _13865_/Y _13878_/D VGND VGND VPWR VPWR _13879_/B sky130_fd_sc_hd__or4_4
XFILLER_35_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16060__B1 _11545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15617_ _15740_/A VGND VGND VPWR VPWR _15617_/X sky130_fd_sc_hd__buf_2
X_18405_ _16459_/Y _23819_/Q _16467_/Y _23816_/Q VGND VGND VPWR VPWR _18405_/X sky130_fd_sc_hd__a2bb2o_4
X_12829_ _22377_/A VGND VGND VPWR VPWR _12829_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16597_ _16234_/A VGND VGND VPWR VPWR _16597_/X sky130_fd_sc_hd__buf_2
X_19385_ _19385_/A VGND VGND VPWR VPWR _19385_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15548_ _19825_/A VGND VGND VPWR VPWR _19452_/A sky130_fd_sc_hd__buf_2
X_18336_ _18299_/B _18258_/X _18237_/X _18333_/Y VGND VGND VPWR VPWR _18336_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22684__A1 _22539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23740__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18267_ _23866_/Q _18266_/Y VGND VGND VPWR VPWR _18267_/X sky130_fd_sc_hd__or2_4
X_15479_ HWDATA[25] VGND VGND VPWR VPWR _15479_/X sky130_fd_sc_hd__buf_2
X_17218_ _17217_/Y _17213_/X _16556_/X _17213_/A VGND VGND VPWR VPWR _24012_/D sky130_fd_sc_hd__a2bb2o_4
X_18198_ _23871_/Q VGND VGND VPWR VPWR _18198_/Y sky130_fd_sc_hd__inv_2
X_17149_ _17129_/A _17145_/X _17148_/Y VGND VGND VPWR VPWR _24035_/D sky130_fd_sc_hd__and3_4
XANTENNA__24946__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20160_ _20192_/B VGND VGND VPWR VPWR _20160_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15469__A3 _15468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21538__C _21538_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15874__B1 _11585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22739__A2 _21576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13618__A _13618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20091_ _23095_/Q VGND VGND VPWR VPWR _21142_/B sky130_fd_sc_hd__inv_2
XANTENNA__19065__B1 _19041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12688__B1 _12666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12522__A _12408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18812__B1 _18740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14753__A1_N _24699_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15626__B1 _15386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23850_ _23845_/CLK _23850_/D HRESETn VGND VGND VPWR VPWR _18322_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22801_ _22777_/Y _22781_/X _22785_/X _22801_/D VGND VGND VPWR VPWR HRDATA[24] sky130_fd_sc_hd__or4_4
XFILLER_77_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23781_ _25183_/CLK _23781_/D HRESETn VGND VGND VPWR VPWR RsTx_S1 sky130_fd_sc_hd__dfstp_4
X_20993_ _20998_/A _20993_/B VGND VGND VPWR VPWR _20993_/X sky130_fd_sc_hd__or2_4
XANTENNA__23899__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22732_ _16162_/A _22953_/B VGND VGND VPWR VPWR _22732_/X sky130_fd_sc_hd__and2_4
XFILLER_129_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20922__A1 _20413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23828__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20922__B2 _21638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21570__A _21570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22663_ _12617_/Y _20910_/X _12851_/Y _22029_/X VGND VGND VPWR VPWR _22663_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22124__B1 _15889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24402_ _24620_/CLK _15891_/X HRESETn VGND VGND VPWR VPWR _15889_/A sky130_fd_sc_hd__dfrtp_4
X_21614_ _21626_/A _21614_/B _21613_/X VGND VGND VPWR VPWR _21614_/X sky130_fd_sc_hd__and3_4
XFILLER_107_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_230_0_HCLK clkbuf_8_231_0_HCLK/A VGND VGND VPWR VPWR _24606_/CLK sky130_fd_sc_hd__clkbuf_1
X_22594_ _21051_/X VGND VGND VPWR VPWR _22597_/A sky130_fd_sc_hd__buf_2
X_24333_ _24333_/CLK _24333_/D HRESETn VGND VGND VPWR VPWR _24333_/Q sky130_fd_sc_hd__dfrtp_4
X_21545_ _11623_/Y _11986_/X _15991_/Y _21544_/X VGND VGND VPWR VPWR _21545_/X sky130_fd_sc_hd__o22a_4
XFILLER_21_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11601__A HWDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24264_ _24264_/CLK _16281_/X HRESETn VGND VGND VPWR VPWR _24264_/Q sky130_fd_sc_hd__dfrtp_4
X_21476_ _21155_/A _21474_/X _21475_/X VGND VGND VPWR VPWR _21476_/X sky130_fd_sc_hd__and3_4
XFILLER_5_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20914__A _21591_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17495__A _22473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23215_ _23293_/CLK _23215_/D VGND VGND VPWR VPWR _19776_/A sky130_fd_sc_hd__dfxtp_4
X_20427_ _21285_/A _20416_/X _20425_/X _20426_/X VGND VGND VPWR VPWR _20428_/A sky130_fd_sc_hd__o22a_4
XANTENNA__21729__B _20832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24687__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24195_ _24192_/CLK _24195_/D HRESETn VGND VGND VPWR VPWR _16462_/A sky130_fd_sc_hd__dfrtp_4
X_23146_ _25067_/CLK _23146_/D VGND VGND VPWR VPWR _23146_/Q sky130_fd_sc_hd__dfxtp_4
X_20358_ _20357_/X VGND VGND VPWR VPWR _20358_/X sky130_fd_sc_hd__buf_2
XFILLER_122_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24616__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15865__B1 _15777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20289_ _20289_/A _20288_/Y _20278_/X VGND VGND VPWR VPWR _20289_/X sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_4_2_0_HCLK_A clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23077_ _23624_/CLK _20132_/X VGND VGND VPWR VPWR _23077_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_136_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22028_ _22028_/A _22025_/X _22026_/X _22027_/X VGND VGND VPWR VPWR _22028_/X sky130_fd_sc_hd__or4_4
XFILLER_0_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22532__A2_N _22530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14850_ _24149_/Q VGND VGND VPWR VPWR _14850_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15743__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13801_ _13869_/A VGND VGND VPWR VPWR _13866_/A sky130_fd_sc_hd__inv_2
XFILLER_5_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15632__A3 _15522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14781_ _24115_/Q VGND VGND VPWR VPWR _14781_/Y sky130_fd_sc_hd__inv_2
X_11993_ _11992_/Y _11990_/X _11607_/X _11990_/X VGND VGND VPWR VPWR _11993_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23979_ _23979_/CLK _17443_/X HRESETn VGND VGND VPWR VPWR _23979_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16520_ _16520_/A VGND VGND VPWR VPWR _16520_/Y sky130_fd_sc_hd__inv_2
X_13732_ _13732_/A _13732_/B _13730_/X _13732_/D VGND VGND VPWR VPWR _13735_/A sky130_fd_sc_hd__and4_4
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11654__B2 _23922_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22576__A _22576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20913__B2 _20827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_40_0_HCLK clkbuf_6_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_40_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_16451_ HWDATA[9] VGND VGND VPWR VPWR _16451_/X sky130_fd_sc_hd__buf_2
X_13663_ _13663_/A VGND VGND VPWR VPWR _13663_/X sky130_fd_sc_hd__buf_2
XFILLER_73_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22115__B1 _21062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15402_ _21285_/A _15396_/X _15286_/X _15401_/X VGND VGND VPWR VPWR _24586_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20808__B _13618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12614_ _25041_/Q VGND VGND VPWR VPWR _12737_/A sky130_fd_sc_hd__inv_2
X_19170_ _18763_/X VGND VGND VPWR VPWR _19170_/X sky130_fd_sc_hd__buf_2
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16382_ _16381_/Y _16379_/X _16211_/X _16379_/X VGND VGND VPWR VPWR _24225_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22666__A1 _12854_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13594_ _13580_/A VGND VGND VPWR VPWR _13594_/X sky130_fd_sc_hd__buf_2
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18121_ _21586_/B _18118_/X _23881_/Q _18118_/X VGND VGND VPWR VPWR _23882_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15333_ _15353_/A VGND VGND VPWR VPWR _15333_/X sky130_fd_sc_hd__buf_2
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12545_ _12544_/Y _24533_/Q _12544_/Y _24533_/Q VGND VGND VPWR VPWR _12545_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14094__A _13398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12607__A _25054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18052_ _17631_/Y _18034_/X _17636_/A _18035_/Y VGND VGND VPWR VPWR _18052_/X sky130_fd_sc_hd__o22a_4
X_15264_ _23766_/Q _15260_/X _15251_/Y _13730_/X _15262_/X VGND VGND VPWR VPWR _15264_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_32_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12476_ _12412_/C _12480_/B _12475_/Y VGND VGND VPWR VPWR _12476_/X sky130_fd_sc_hd__o21a_4
X_17003_ _16181_/Y _24042_/Q _16181_/Y _24042_/Q VGND VGND VPWR VPWR _17003_/X sky130_fd_sc_hd__a2bb2o_4
X_14215_ _21073_/A VGND VGND VPWR VPWR _14215_/Y sky130_fd_sc_hd__inv_2
X_15195_ _14903_/Y _15159_/A VGND VGND VPWR VPWR _15229_/A sky130_fd_sc_hd__or2_4
XFILLER_126_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14146_ _24839_/Q _12051_/X _14145_/X VGND VGND VPWR VPWR _14147_/A sky130_fd_sc_hd__a21o_4
XFILLER_10_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24357__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14541__B _14437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15856__B1 _15855_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19047__B1 _18932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14077_ _14077_/A VGND VGND VPWR VPWR _14077_/Y sky130_fd_sc_hd__inv_2
X_18954_ _18952_/Y _18950_/X _18953_/X _18950_/X VGND VGND VPWR VPWR _23507_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17058__C1 _17057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13028_ _13045_/A _13028_/B VGND VGND VPWR VPWR _13028_/X sky130_fd_sc_hd__or2_4
X_17905_ _17969_/A _17905_/B _17904_/X VGND VGND VPWR VPWR _17905_/X sky130_fd_sc_hd__or3_4
X_18885_ _18882_/Y _18877_/X _18883_/X _18884_/X VGND VGND VPWR VPWR _23532_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15608__B1 _11566_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17836_ _17732_/A VGND VGND VPWR VPWR _17968_/A sky130_fd_sc_hd__buf_2
XFILLER_39_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_122_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_245_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__19784__A1_N _19783_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16281__B1 _15978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17767_ _17767_/A VGND VGND VPWR VPWR _17767_/X sky130_fd_sc_hd__buf_2
XFILLER_81_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14979_ _24713_/Q _14979_/B VGND VGND VPWR VPWR _14981_/B sky130_fd_sc_hd__or2_4
XANTENNA__18964__A _18711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23992__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19506_ _19859_/A VGND VGND VPWR VPWR _19506_/X sky130_fd_sc_hd__buf_2
X_16718_ _16718_/A VGND VGND VPWR VPWR _17558_/B sky130_fd_sc_hd__inv_2
X_17698_ _17698_/A _23430_/Q VGND VGND VPWR VPWR _17699_/C sky130_fd_sc_hd__or2_4
XANTENNA__23921__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20904__B2 _20827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21390__A _21235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25145__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19437_ _19436_/Y _19432_/X _19392_/X _19417_/Y VGND VGND VPWR VPWR _19437_/X sky130_fd_sc_hd__a2bb2o_4
X_16649_ _16649_/A VGND VGND VPWR VPWR _16649_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19368_ _13306_/B VGND VGND VPWR VPWR _19368_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20668__B1 _24184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18319_ _18262_/A VGND VGND VPWR VPWR _18319_/X sky130_fd_sc_hd__buf_2
XANTENNA__13620__B _13619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19299_ _19298_/Y _19296_/X _11860_/X _19296_/X VGND VGND VPWR VPWR _19299_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22933__B _22933_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14435__C _14369_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21330_ _21350_/A _21328_/X _21330_/C VGND VGND VPWR VPWR _21330_/X sky130_fd_sc_hd__and3_4
XANTENNA__20683__A3 _13543_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_60_0_HCLK clkbuf_7_30_0_HCLK/X VGND VGND VPWR VPWR _23969_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16931__B _16927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21261_ _21247_/Y _21259_/Y _21793_/A VGND VGND VPWR VPWR _21261_/X sky130_fd_sc_hd__o21a_4
XFILLER_102_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15828__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24780__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21549__B _16042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14732__A _14732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23811__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23000_ _15463_/X _22999_/X _22251_/X _24426_/Q _15824_/A VGND VGND VPWR VPWR _23001_/B
+ sky130_fd_sc_hd__a32o_4
X_20212_ _15260_/A _20212_/B _23771_/Q _20212_/D VGND VGND VPWR VPWR _20266_/A sky130_fd_sc_hd__and4_4
XFILLER_132_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21192_ _22045_/B VGND VGND VPWR VPWR _21192_/X sky130_fd_sc_hd__buf_2
XANTENNA__24098__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20143_ _23073_/Q VGND VGND VPWR VPWR _20143_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24027__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20074_ _20074_/A VGND VGND VPWR VPWR _22084_/B sky130_fd_sc_hd__inv_2
X_24951_ _24957_/CLK _24951_/D HRESETn VGND VGND VPWR VPWR _11650_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_131_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16659__A _16643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15563__A _15556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23902_ _23353_/CLK _23902_/D HRESETn VGND VGND VPWR VPWR _18023_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24882_ _24884_/CLK _14003_/Y HRESETn VGND VGND VPWR VPWR _13925_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16272__B1 _22477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15614__A3 _15497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23833_ _23828_/CLK _23833_/D HRESETn VGND VGND VPWR VPWR _23833_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22345__B1 _21886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23764_ _24644_/CLK _20263_/X HRESETn VGND VGND VPWR VPWR _23764_/Q sky130_fd_sc_hd__dfrtp_4
X_20976_ _21130_/A VGND VGND VPWR VPWR _20980_/A sky130_fd_sc_hd__buf_2
XANTENNA__23662__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_27_0_HCLK clkbuf_5_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22715_ _20512_/Y _22610_/X _23748_/Q _22657_/X VGND VGND VPWR VPWR _22715_/X sky130_fd_sc_hd__a2bb2o_4
X_23695_ _24161_/CLK _20421_/Y HRESETn VGND VGND VPWR VPWR _21020_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_41_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14907__A _24274_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22646_ _22646_/A VGND VGND VPWR VPWR _22646_/X sky130_fd_sc_hd__buf_2
XANTENNA__21320__A1 _12534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22577_ _24273_/Q _22477_/B _22338_/X VGND VGND VPWR VPWR _22577_/X sky130_fd_sc_hd__o21a_4
X_12330_ _12328_/A _12329_/A _12328_/Y _12329_/Y VGND VGND VPWR VPWR _12337_/B sky130_fd_sc_hd__o22a_4
X_24316_ _24055_/CLK _24316_/D HRESETn VGND VGND VPWR VPWR _24316_/Q sky130_fd_sc_hd__dfrtp_4
X_21528_ _21396_/A _21528_/B _21528_/C VGND VGND VPWR VPWR _21528_/X sky130_fd_sc_hd__or3_4
X_12261_ _12261_/A _12261_/B _12260_/X VGND VGND VPWR VPWR _12261_/X sky130_fd_sc_hd__and3_4
XANTENNA__15738__A _15418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24247_ _24213_/CLK _16324_/X HRESETn VGND VGND VPWR VPWR _24247_/Q sky130_fd_sc_hd__dfrtp_4
X_21459_ _21348_/A _21459_/B VGND VGND VPWR VPWR _21459_/X sky130_fd_sc_hd__or2_4
XFILLER_5_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14000_ _13925_/B _14000_/B VGND VGND VPWR VPWR _14000_/Y sky130_fd_sc_hd__nor2_4
XFILLER_123_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24450__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12192_ _12192_/A _12192_/B VGND VGND VPWR VPWR _12193_/B sky130_fd_sc_hd__or2_4
XFILLER_135_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15457__B _15456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24178_ _24177_/CLK _24178_/D HRESETn VGND VGND VPWR VPWR _16505_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15838__B1 _15837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23129_ _23993_/CLK _20004_/X VGND VGND VPWR VPWR _23129_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_110_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21475__A _21342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15951_ _15950_/Y _15948_/X _15770_/X _15948_/X VGND VGND VPWR VPWR _24380_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14902_ _24671_/Q _14900_/Y _24677_/Q _14901_/Y VGND VGND VPWR VPWR _14905_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15882_ _24405_/Q VGND VGND VPWR VPWR _15882_/Y sky130_fd_sc_hd__inv_2
X_18670_ _18670_/A VGND VGND VPWR VPWR _18670_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16263__B1 _16261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17621_ _17619_/A _17615_/B _17620_/Y VGND VGND VPWR VPWR _17621_/X sky130_fd_sc_hd__and3_4
X_14833_ _24146_/Q VGND VGND VPWR VPWR _14833_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14813__A1 _24698_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11506__A _23763_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14764_ _15019_/A _16655_/A _15019_/A _16655_/A VGND VGND VPWR VPWR _14764_/X sky130_fd_sc_hd__a2bb2o_4
X_17552_ _17554_/B VGND VGND VPWR VPWR _17553_/B sky130_fd_sc_hd__inv_2
XANTENNA__22887__A1 _22931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11976_ _11975_/Y _11971_/X _11631_/X _11971_/X VGND VGND VPWR VPWR _11976_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20819__A _20818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13715_ _24649_/Q VGND VGND VPWR VPWR _13770_/A sky130_fd_sc_hd__buf_2
X_16503_ _24179_/Q VGND VGND VPWR VPWR _22695_/A sky130_fd_sc_hd__inv_2
XANTENNA__20898__B1 _20897_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17483_ _17483_/A _16702_/Y VGND VGND VPWR VPWR _17502_/C sky130_fd_sc_hd__or2_4
XANTENNA__15920__B _15919_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14695_ _14869_/A VGND VGND VPWR VPWR _15064_/A sky130_fd_sc_hd__buf_2
X_19222_ _19220_/Y _19218_/X _19221_/X _19218_/X VGND VGND VPWR VPWR _23411_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13646_ _13643_/Y _13639_/X _13645_/X _13639_/X VGND VGND VPWR VPWR _24941_/D sky130_fd_sc_hd__a2bb2o_4
X_16434_ _16452_/A VGND VGND VPWR VPWR _16434_/X sky130_fd_sc_hd__buf_2
XFILLER_34_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16365_ _16363_/Y _16359_/X _15978_/X _16364_/X VGND VGND VPWR VPWR _16365_/X sky130_fd_sc_hd__a2bb2o_4
X_19153_ _19153_/A VGND VGND VPWR VPWR _19153_/X sky130_fd_sc_hd__buf_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13577_ _13572_/X _13553_/X _13575_/Y _13576_/X _13566_/C VGND VGND VPWR VPWR _24960_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22753__B _22587_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21311__B2 _20759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15316_ _15315_/X VGND VGND VPWR VPWR _21019_/A sky130_fd_sc_hd__buf_2
X_18104_ _18104_/A _18104_/B VGND VGND VPWR VPWR _18104_/Y sky130_fd_sc_hd__nor2_4
X_12528_ _12527_/X VGND VGND VPWR VPWR _12528_/Y sky130_fd_sc_hd__inv_2
X_16296_ _16296_/A VGND VGND VPWR VPWR _16296_/Y sky130_fd_sc_hd__inv_2
X_19084_ _19078_/Y VGND VGND VPWR VPWR _19084_/X sky130_fd_sc_hd__buf_2
XFILLER_9_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24538__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_47_0_HCLK clkbuf_7_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_95_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15247_ _15260_/A VGND VGND VPWR VPWR _15247_/X sky130_fd_sc_hd__buf_2
X_18035_ _18034_/X VGND VGND VPWR VPWR _18035_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15648__A _15418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12459_ _25093_/Q _12458_/Y VGND VGND VPWR VPWR _12459_/X sky130_fd_sc_hd__or2_4
XANTENNA__13001__B1 _12896_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15178_ _15165_/A _15178_/B _15177_/Y VGND VGND VPWR VPWR _24667_/D sky130_fd_sc_hd__and3_4
XANTENNA__22811__A1 _21561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24191__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18959__A _16291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15829__B1 _15828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12760__C1 _12674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14129_ _14126_/X _14128_/Y _13332_/A _14126_/X VGND VGND VPWR VPWR _24848_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24120__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19986_ _23135_/Q VGND VGND VPWR VPWR _19986_/Y sky130_fd_sc_hd__inv_2
X_18937_ _23512_/Q VGND VGND VPWR VPWR _18937_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18868_ _13259_/B VGND VGND VPWR VPWR _18868_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17819_ _17781_/A _23419_/Q VGND VGND VPWR VPWR _17819_/X sky130_fd_sc_hd__or2_4
X_18799_ _18797_/Y _18798_/X _18706_/X _18798_/X VGND VGND VPWR VPWR _18799_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14804__B2 _24153_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22928__B _23020_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20830_ _21716_/B _20828_/X _24461_/Q _22859_/A VGND VGND VPWR VPWR _20830_/X sky130_fd_sc_hd__o22a_4
XFILLER_39_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20761_ _21448_/B VGND VGND VPWR VPWR _22014_/B sky130_fd_sc_hd__buf_2
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16557__B2 _16493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21550__B2 _21107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22500_ _22500_/A _22499_/X VGND VGND VPWR VPWR _22500_/Y sky130_fd_sc_hd__nor2_4
XFILLER_56_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23480_ _23479_/CLK _19028_/X VGND VGND VPWR VPWR _19027_/A sky130_fd_sc_hd__dfxtp_4
X_20692_ _11914_/X _20691_/B VGND VGND VPWR VPWR _20692_/X sky130_fd_sc_hd__and2_4
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22431_ _16183_/A _22505_/A VGND VGND VPWR VPWR _22431_/X sky130_fd_sc_hd__and2_4
XANTENNA__24961__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25150_ _24824_/CLK _25150_/D HRESETn VGND VGND VPWR VPWR _25150_/Q sky130_fd_sc_hd__dfrtp_4
X_22362_ _22116_/X _22361_/X _21974_/X _25202_/Q _22118_/X VGND VGND VPWR VPWR _22362_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24279__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24101_ _24101_/CLK _16664_/X HRESETn VGND VGND VPWR VPWR _14726_/A sky130_fd_sc_hd__dfrtp_4
X_21313_ _21308_/X _21312_/X VGND VGND VPWR VPWR _21323_/C sky130_fd_sc_hd__and2_4
XFILLER_136_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24208__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25081_ _25097_/CLK _25081_/D HRESETn VGND VGND VPWR VPWR _25081_/Q sky130_fd_sc_hd__dfrtp_4
X_22293_ _22254_/X _22262_/X _22270_/Y _22292_/X VGND VGND VPWR VPWR HRDATA[10] sky130_fd_sc_hd__a211o_4
XANTENNA__15532__A2 _15319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24032_ _24055_/CLK _17156_/X HRESETn VGND VGND VPWR VPWR _24032_/Q sky130_fd_sc_hd__dfrtp_4
X_21244_ _21396_/A _21244_/B _21243_/X VGND VGND VPWR VPWR _21244_/X sky130_fd_sc_hd__or3_4
XFILLER_11_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_4_0_HCLK clkbuf_6_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_4_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21175_ _20777_/X VGND VGND VPWR VPWR _21175_/X sky130_fd_sc_hd__buf_2
XFILLER_78_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20126_ _17982_/A _20119_/X _19808_/X _23080_/Q _20117_/X VGND VGND VPWR VPWR _23080_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22566__B1 _20800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20057_ _20054_/X _15410_/X _13665_/A _21649_/B _20055_/X VGND VGND VPWR VPWR _23108_/D
+ sky130_fd_sc_hd__a32o_4
X_24934_ _24974_/CLK _24934_/D HRESETn VGND VGND VPWR VPWR _24934_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23843__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16245__B1 _15837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25067__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24865_ _24870_/CLK _14063_/X HRESETn VGND VGND VPWR VPWR _14062_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__22838__B _23008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11830_ _11830_/A VGND VGND VPWR VPWR _11830_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23816_ _23824_/CLK _18554_/X HRESETn VGND VGND VPWR VPWR _23816_/Q sky130_fd_sc_hd__dfrtp_4
X_24796_ _24859_/CLK _14276_/X HRESETn VGND VGND VPWR VPWR _24796_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23015__A _22982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11761_/A _11761_/B VGND VGND VPWR VPWR _11761_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__19212__B _16127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23747_ _24177_/CLK _23747_/D HRESETn VGND VGND VPWR VPWR _13524_/B sky130_fd_sc_hd__dfrtp_4
X_20959_ _17646_/A VGND VGND VPWR VPWR _20965_/A sky130_fd_sc_hd__buf_2
XFILLER_57_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13498_/Y _13499_/Y VGND VGND VPWR VPWR _13500_/X sky130_fd_sc_hd__and2_4
XPHY_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14480_/A VGND VGND VPWR VPWR _14480_/X sky130_fd_sc_hd__buf_2
XFILLER_42_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _13566_/C _23923_/Q _13572_/A _11691_/Y VGND VGND VPWR VPWR _11692_/X sky130_fd_sc_hd__o22a_4
XPHY_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23678_ _24728_/CLK _20396_/X HRESETn VGND VGND VPWR VPWR _23678_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _24935_/Q VGND VGND VPWR VPWR _22271_/A sky130_fd_sc_hd__inv_2
XPHY_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22629_ _22629_/A VGND VGND VPWR VPWR _22629_/X sky130_fd_sc_hd__buf_2
XPHY_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16150_ _16149_/Y _16145_/X _15756_/X _16145_/X VGND VGND VPWR VPWR _24316_/D sky130_fd_sc_hd__a2bb2o_4
X_13362_ _13362_/A _13328_/X VGND VGND VPWR VPWR _13363_/A sky130_fd_sc_hd__nor2_4
XFILLER_10_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15101_ _24678_/Q VGND VGND VPWR VPWR _15129_/A sky130_fd_sc_hd__inv_2
X_12313_ _12313_/A VGND VGND VPWR VPWR _12412_/D sky130_fd_sc_hd__inv_2
X_16081_ _16080_/Y _16076_/X _15777_/X _16076_/X VGND VGND VPWR VPWR _16081_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15468__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13293_ _13261_/A _18986_/A VGND VGND VPWR VPWR _13293_/X sky130_fd_sc_hd__or2_4
X_15032_ _14736_/X _15036_/B _15031_/Y VGND VGND VPWR VPWR _24701_/D sky130_fd_sc_hd__o21a_4
X_12244_ _12174_/A _12244_/B VGND VGND VPWR VPWR _12245_/C sky130_fd_sc_hd__nand2_4
XFILLER_107_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19840_ _19862_/A _14541_/X VGND VGND VPWR VPWR _19841_/A sky130_fd_sc_hd__and2_4
X_12175_ _12175_/A _12149_/Y _12175_/C VGND VGND VPWR VPWR _12183_/A sky130_fd_sc_hd__or3_4
XFILLER_122_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16484__B1 _16243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19771_ _23217_/Q VGND VGND VPWR VPWR _21329_/B sky130_fd_sc_hd__inv_2
X_16983_ _24308_/Q _24046_/Q _16169_/Y _16982_/Y VGND VGND VPWR VPWR _16990_/A sky130_fd_sc_hd__o22a_4
X_18722_ _18721_/Y _18719_/X _18700_/X _18719_/X VGND VGND VPWR VPWR _18722_/X sky130_fd_sc_hd__a2bb2o_4
X_15934_ _15933_/Y _15929_/X _15756_/X _15929_/X VGND VGND VPWR VPWR _24387_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19422__B1 _19421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21933__A _20980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18653_ _18652_/Y _18650_/X _15554_/X _18650_/X VGND VGND VPWR VPWR _18653_/X sky130_fd_sc_hd__a2bb2o_4
X_15865_ _15864_/Y _15860_/X _15777_/X _15860_/X VGND VGND VPWR VPWR _15865_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17984__B1 _22450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17604_ _17595_/C _17607_/B VGND VGND VPWR VPWR _17605_/C sky130_fd_sc_hd__nand2_4
X_14816_ _24133_/Q VGND VGND VPWR VPWR _14816_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18584_ _16343_/Y _18503_/A _24243_/Q _18491_/A VGND VGND VPWR VPWR _18587_/B sky130_fd_sc_hd__a2bb2o_4
X_15796_ _12827_/Y _15795_/X _15393_/X _15795_/X VGND VGND VPWR VPWR _24434_/D sky130_fd_sc_hd__a2bb2o_4
X_17535_ _17535_/A VGND VGND VPWR VPWR _17535_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15650__B _15459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11959_ _25155_/Q VGND VGND VPWR VPWR _11959_/Y sky130_fd_sc_hd__inv_2
X_14747_ _14747_/A VGND VGND VPWR VPWR _14747_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21532__B2 _22548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_10_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_14678_ _14677_/X VGND VGND VPWR VPWR _14678_/Y sky130_fd_sc_hd__inv_2
X_17466_ _17466_/A VGND VGND VPWR VPWR _21805_/A sky130_fd_sc_hd__inv_2
XFILLER_127_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24719__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19205_ _19203_/Y _19204_/X _19115_/X _19204_/X VGND VGND VPWR VPWR _19205_/X sky130_fd_sc_hd__a2bb2o_4
X_13629_ _16042_/A VGND VGND VPWR VPWR _22314_/B sky130_fd_sc_hd__buf_2
X_16417_ _16416_/Y _16414_/X _15484_/X _16414_/X VGND VGND VPWR VPWR _16417_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17397_ _17396_/X VGND VGND VPWR VPWR _23992_/D sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_5_5_0_HCLK_A clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12067__A _11956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20099__B2 _20098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19136_ _19136_/A VGND VGND VPWR VPWR _19136_/Y sky130_fd_sc_hd__inv_2
X_16348_ _16345_/Y _16347_/X _16179_/X _16347_/X VGND VGND VPWR VPWR _16348_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24372__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16279_ HWDATA[10] VGND VGND VPWR VPWR _16279_/X sky130_fd_sc_hd__buf_2
X_19067_ _19066_/Y _19064_/X _18953_/X _19064_/X VGND VGND VPWR VPWR _19067_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24301__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16711__B2 _16710_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21048__B1 _25191_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18018_ _23903_/Q VGND VGND VPWR VPWR _18018_/X sky130_fd_sc_hd__buf_2
XFILLER_12_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22378__A2_N _22259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12733__C1 _12666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22796__B1 _12332_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18689__A _23598_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_134_0_HCLK clkbuf_7_67_0_HCLK/X VGND VGND VPWR VPWR _23416_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_8_197_0_HCLK clkbuf_7_98_0_HCLK/X VGND VGND VPWR VPWR _24162_/CLK sky130_fd_sc_hd__clkbuf_1
X_19969_ _19969_/A VGND VGND VPWR VPWR _19982_/A sky130_fd_sc_hd__inv_2
XFILLER_41_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22980_ _22980_/A _22418_/X VGND VGND VPWR VPWR _22980_/X sky130_fd_sc_hd__and2_4
XFILLER_95_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25160__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21931_ _21340_/A _21931_/B VGND VGND VPWR VPWR _21933_/B sky130_fd_sc_hd__or2_4
XANTENNA__21843__A _20782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24650_ _24654_/CLK _24650_/D HRESETn VGND VGND VPWR VPWR _24650_/Q sky130_fd_sc_hd__dfrtp_4
X_21862_ _21715_/X _21859_/X _22547_/A _21861_/X VGND VGND VPWR VPWR _21863_/A sky130_fd_sc_hd__o22a_4
XANTENNA__16673__A1_N _14754_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13056__A3 _13054_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23601_ _23992_/CLK _18683_/X VGND VGND VPWR VPWR _23601_/Q sky130_fd_sc_hd__dfxtp_4
X_20813_ _15455_/X VGND VGND VPWR VPWR _21565_/A sky130_fd_sc_hd__inv_2
XFILLER_93_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24581_ _24017_/CLK _15434_/X HRESETn VGND VGND VPWR VPWR _13546_/A sky130_fd_sc_hd__dfrtp_4
X_21793_ _21793_/A _21792_/X VGND VGND VPWR VPWR _21857_/C sky130_fd_sc_hd__and2_4
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13361__A _22745_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23532_ _23531_/CLK _23532_/D VGND VGND VPWR VPWR _18882_/A sky130_fd_sc_hd__dfxtp_4
X_20744_ _20800_/A VGND VGND VPWR VPWR _20744_/X sky130_fd_sc_hd__buf_2
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23463_ _23419_/CLK _23463_/D VGND VGND VPWR VPWR _19075_/A sky130_fd_sc_hd__dfxtp_4
X_20675_ _23756_/Q VGND VGND VPWR VPWR _20675_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25202_ _23969_/CLK _11595_/X HRESETn VGND VGND VPWR VPWR _25202_/Q sky130_fd_sc_hd__dfrtp_4
X_22414_ _22175_/A _22412_/Y _22349_/B _22413_/X VGND VGND VPWR VPWR _22414_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12408__C _12408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23394_ _23411_/CLK _19272_/X VGND VGND VPWR VPWR _23394_/Q sky130_fd_sc_hd__dfxtp_4
X_25133_ _25084_/CLK _12190_/X HRESETn VGND VGND VPWR VPWR _25133_/Q sky130_fd_sc_hd__dfrtp_4
X_22345_ _22280_/X _22343_/X _21886_/X _22344_/X VGND VGND VPWR VPWR _22345_/X sky130_fd_sc_hd__o22a_4
XFILLER_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23028__A1 _22429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24042__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16611__A1_N _14836_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_30_0_HCLK clkbuf_7_30_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_30_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_25064_ _25061_/CLK _25064_/D HRESETn VGND VGND VPWR VPWR _12547_/A sky130_fd_sc_hd__dfrtp_4
X_22276_ _22275_/X VGND VGND VPWR VPWR _22512_/A sky130_fd_sc_hd__inv_2
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_93_0_HCLK clkbuf_6_46_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_93_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_24015_ _24017_/CLK _17211_/X HRESETn VGND VGND VPWR VPWR _24015_/Q sky130_fd_sc_hd__dfrtp_4
X_21227_ _21227_/A _19525_/Y VGND VGND VPWR VPWR _21227_/X sky130_fd_sc_hd__or2_4
XANTENNA__14951__A2_N _22477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15269__A1 _14100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16466__B1 _15992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21158_ _21158_/A _21158_/B VGND VGND VPWR VPWR _21160_/B sky130_fd_sc_hd__or2_4
XFILLER_78_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20109_ _23088_/Q VGND VGND VPWR VPWR _20109_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13536__A _23742_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13980_ _24887_/Q _13941_/X _24887_/Q _13941_/X VGND VGND VPWR VPWR _13981_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22003__A2 _21976_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21089_ _17215_/Y _21043_/X _23656_/Q _21088_/X VGND VGND VPWR VPWR _21090_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12440__A _12417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12931_ _12922_/A _12931_/B _12930_/X VGND VGND VPWR VPWR _12932_/A sky130_fd_sc_hd__or3_4
XFILLER_92_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24917_ _24923_/CLK _13703_/X HRESETn VGND VGND VPWR VPWR _24917_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12862_ _22921_/A _12849_/Y _12972_/A _15797_/A VGND VGND VPWR VPWR _12865_/C sky130_fd_sc_hd__a2bb2o_4
X_15650_ _11944_/X _15459_/A VGND VGND VPWR VPWR _15650_/X sky130_fd_sc_hd__or2_4
XFILLER_46_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24848_ _24847_/CLK _24848_/D HRESETn VGND VGND VPWR VPWR MSO_S2 sky130_fd_sc_hd__dfrtp_4
X_11813_ _11777_/X _11823_/A _11817_/B VGND VGND VPWR VPWR _11818_/A sky130_fd_sc_hd__o21a_4
X_14601_ _24732_/Q VGND VGND VPWR VPWR _19946_/C sky130_fd_sc_hd__buf_2
X_15581_ _15740_/A VGND VGND VPWR VPWR _15582_/A sky130_fd_sc_hd__buf_2
X_12793_ _25005_/Q VGND VGND VPWR VPWR _12793_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24883__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24779_ _23618_/CLK _24779_/D HRESETn VGND VGND VPWR VPWR _20331_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14367__A HREADY VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__A _13271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14441_/A VGND VGND VPWR VPWR _20994_/A sky130_fd_sc_hd__inv_2
X_17320_ _17320_/A _17264_/Y _17319_/Y _17415_/A VGND VGND VPWR VPWR _17324_/B sky130_fd_sc_hd__or4_4
XPHY_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _18065_/C _18085_/A _18065_/C _18085_/A VGND VGND VPWR VPWR _11745_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14462_/X VGND VGND VPWR VPWR _14463_/Y sky130_fd_sc_hd__inv_2
X_17251_ _17251_/A VGND VGND VPWR VPWR _17251_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ _11673_/A _23920_/Q _11673_/Y _22272_/A VGND VGND VPWR VPWR _11682_/B sky130_fd_sc_hd__o22a_4
XPHY_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13414_ _24931_/Q _13413_/Y _13408_/Y _14377_/A VGND VGND VPWR VPWR _13414_/X sky130_fd_sc_hd__a2bb2o_4
X_16202_ _16202_/A VGND VGND VPWR VPWR _16202_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21278__B1 _20807_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17182_ _23678_/Q _17182_/B VGND VGND VPWR VPWR _20394_/A sky130_fd_sc_hd__or2_4
XFILLER_35_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14394_ _14394_/A _14393_/Y VGND VGND VPWR VPWR _14394_/X sky130_fd_sc_hd__or2_4
XFILLER_31_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18143__B1 _16056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16133_ _22999_/A VGND VGND VPWR VPWR _16133_/Y sky130_fd_sc_hd__inv_2
X_13345_ _13343_/Y _13339_/X _11620_/X _13344_/X VGND VGND VPWR VPWR _24992_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16064_ _16071_/A VGND VGND VPWR VPWR _16064_/X sky130_fd_sc_hd__buf_2
XANTENNA__14704__B1 _14703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13276_ _13182_/A _19051_/A VGND VGND VPWR VPWR _13276_/X sky130_fd_sc_hd__or2_4
XANTENNA__20832__A _20832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15015_ _15003_/B _14982_/X _15003_/A VGND VGND VPWR VPWR _15015_/X sky130_fd_sc_hd__o21a_4
X_12227_ _12165_/X VGND VGND VPWR VPWR _12227_/X sky130_fd_sc_hd__buf_2
XANTENNA__23765__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_207_0_HCLK clkbuf_8_207_0_HCLK/A VGND VGND VPWR VPWR _24259_/CLK sky130_fd_sc_hd__clkbuf_1
X_19823_ _21781_/B _19814_/X _19821_/X _19822_/X VGND VGND VPWR VPWR _23196_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20104__A2_N _20098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12158_ _12152_/Y VGND VGND VPWR VPWR _12265_/A sky130_fd_sc_hd__buf_2
XANTENNA__15645__B _16127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19754_ _23223_/Q VGND VGND VPWR VPWR _20974_/B sky130_fd_sc_hd__inv_2
XFILLER_68_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12089_ _12089_/A VGND VGND VPWR VPWR _12089_/Y sky130_fd_sc_hd__inv_2
X_16966_ _16966_/A VGND VGND VPWR VPWR _16966_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16209__B1 _15992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22759__A _22681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18705_ _18697_/A VGND VGND VPWR VPWR _18705_/X sky130_fd_sc_hd__buf_2
X_15917_ _11535_/X _15915_/X _15912_/X _24392_/Q _15916_/X VGND VGND VPWR VPWR _15917_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_83_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19685_ _19684_/Y _19680_/X _19641_/X _19680_/A VGND VGND VPWR VPWR _19685_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16897_ _16765_/Y _16895_/X _16896_/Y VGND VGND VPWR VPWR _16897_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24801__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18636_ _21188_/A _11708_/A VGND VGND VPWR VPWR _18636_/X sky130_fd_sc_hd__and2_4
X_15848_ _15846_/Y _15842_/X _15761_/X _15847_/X VGND VGND VPWR VPWR _24419_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24864__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18567_ _16323_/Y _18472_/A _16323_/Y _18472_/A VGND VGND VPWR VPWR _18571_/A sky130_fd_sc_hd__a2bb2o_4
X_15779_ _15746_/A VGND VGND VPWR VPWR _15779_/X sky130_fd_sc_hd__buf_2
XANTENNA__13443__B1 _13441_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13181__A _13271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17518_ _16710_/Y _17518_/B VGND VGND VPWR VPWR _17519_/C sky130_fd_sc_hd__or2_4
XANTENNA__24553__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18498_ _18434_/D _18495_/D VGND VGND VPWR VPWR _18502_/A sky130_fd_sc_hd__or2_4
XFILLER_36_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17449_ _17447_/Y _17460_/B VGND VGND VPWR VPWR _17449_/X sky130_fd_sc_hd__or2_4
XANTENNA__17588__A _21839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20460_ _20460_/A VGND VGND VPWR VPWR _20460_/Y sky130_fd_sc_hd__inv_2
X_19119_ _23447_/Q VGND VGND VPWR VPWR _19119_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20391_ _15278_/Y _20343_/Y _20357_/X _20390_/X VGND VGND VPWR VPWR _20391_/X sky130_fd_sc_hd__a211o_4
X_22130_ _24474_/Q _22524_/B VGND VGND VPWR VPWR _22130_/X sky130_fd_sc_hd__or2_4
XFILLER_12_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_17_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__20742__A _11725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22061_ _22064_/A _22061_/B VGND VGND VPWR VPWR _22061_/X sky130_fd_sc_hd__or2_4
XFILLER_82_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15836__A _24423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22233__A2 _22232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21012_ _21012_/A _19901_/Y VGND VGND VPWR VPWR _21012_/X sky130_fd_sc_hd__or2_4
XFILLER_87_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20795__A2 _20780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12139__A2_N _24560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21573__A _24259_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22963_ _22963_/A VGND VGND VPWR VPWR _22964_/C sky130_fd_sc_hd__inv_2
XFILLER_74_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22388__B _22246_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21914_ _20980_/A _21914_/B _21914_/C VGND VGND VPWR VPWR _21914_/X sky130_fd_sc_hd__and3_4
XANTENNA__15571__A _22884_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24702_ _24706_/CLK _15029_/Y HRESETn VGND VGND VPWR VPWR _24702_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22894_ _24387_/Q _22638_/X VGND VGND VPWR VPWR _22894_/X sky130_fd_sc_hd__or2_4
XFILLER_71_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15423__A1 _15421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24633_ _24641_/CLK _24633_/D HRESETn VGND VGND VPWR VPWR _13754_/B sky130_fd_sc_hd__dfrtp_4
X_21845_ _24472_/Q _22036_/A VGND VGND VPWR VPWR _21845_/X sky130_fd_sc_hd__or2_4
XFILLER_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13091__A _11741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11604__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24294__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24564_ _24573_/CLK _15491_/X HRESETn VGND VGND VPWR VPWR _24564_/Q sky130_fd_sc_hd__dfrtp_4
X_21776_ _21771_/X _21775_/X _14523_/A VGND VGND VPWR VPWR _21776_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_58_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11996__B1 _11612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23515_ _23514_/CLK _23515_/D VGND VGND VPWR VPWR _17838_/B sky130_fd_sc_hd__dfxtp_4
X_20727_ _23666_/D VGND VGND VPWR VPWR _20729_/A sky130_fd_sc_hd__inv_2
XANTENNA__17498__A _17498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24223__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24495_ _24604_/CLK _24495_/D HRESETn VGND VGND VPWR VPWR _24495_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23446_ _24735_/CLK _23446_/D VGND VGND VPWR VPWR _23446_/Q sky130_fd_sc_hd__dfxtp_4
X_20658_ _16497_/Y _20552_/X _20583_/X _20657_/X VGND VGND VPWR VPWR _20658_/X sky130_fd_sc_hd__o22a_4
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23377_ _25002_/CLK _23377_/D VGND VGND VPWR VPWR _13245_/B sky130_fd_sc_hd__dfxtp_4
X_20589_ _20589_/A VGND VGND VPWR VPWR _20589_/Y sky130_fd_sc_hd__inv_2
X_13130_ _13204_/A _23604_/Q VGND VGND VPWR VPWR _13130_/X sky130_fd_sc_hd__or2_4
X_25116_ _25106_/CLK _12254_/Y HRESETn VGND VGND VPWR VPWR _12129_/A sky130_fd_sc_hd__dfrtp_4
X_22328_ _16445_/Y _22230_/A _16658_/Y _22017_/X VGND VGND VPWR VPWR _22328_/X sky130_fd_sc_hd__o22a_4
XFILLER_124_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13061_ _13297_/A _13061_/B VGND VGND VPWR VPWR _13061_/X sky130_fd_sc_hd__or2_4
XANTENNA__15746__A _15746_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25047_ _25046_/CLK _12747_/X HRESETn VGND VGND VPWR VPWR _12648_/A sky130_fd_sc_hd__dfrtp_4
X_22259_ _22259_/A VGND VGND VPWR VPWR _22259_/X sky130_fd_sc_hd__buf_2
XFILLER_69_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21467__B _19677_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22208__A2_N _21707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12012_ _12011_/Y _12007_/X _11643_/X _12007_/X VGND VGND VPWR VPWR _12012_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25082__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16820_ _24084_/Q VGND VGND VPWR VPWR _16863_/A sky130_fd_sc_hd__inv_2
XANTENNA__25011__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_180_0_HCLK clkbuf_7_90_0_HCLK/X VGND VGND VPWR VPWR _24445_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_93_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_37_0_HCLK clkbuf_8_37_0_HCLK/A VGND VGND VPWR VPWR _23374_/CLK sky130_fd_sc_hd__clkbuf_1
X_16751_ _15879_/Y _16833_/A _15879_/Y _16833_/A VGND VGND VPWR VPWR _16756_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12476__A1 _12412_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13963_ _13936_/A VGND VGND VPWR VPWR _13963_/X sky130_fd_sc_hd__buf_2
XFILLER_24_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13673__B1 _13638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21735__B2 _21088_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15702_ _15695_/A VGND VGND VPWR VPWR _15702_/X sky130_fd_sc_hd__buf_2
X_12914_ _12914_/A VGND VGND VPWR VPWR _12914_/Y sky130_fd_sc_hd__inv_2
X_19470_ _19470_/A VGND VGND VPWR VPWR _19470_/Y sky130_fd_sc_hd__inv_2
X_13894_ _13828_/D _13892_/X _13884_/X _13828_/C _13893_/X VGND VGND VPWR VPWR _24911_/D
+ sky130_fd_sc_hd__a32o_4
X_16682_ _16681_/X VGND VGND VPWR VPWR _24092_/D sky130_fd_sc_hd__inv_2
X_18421_ _18420_/Y _18421_/B VGND VGND VPWR VPWR _18427_/B sky130_fd_sc_hd__or2_4
XANTENNA__16611__B1 _16373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12845_ _12845_/A VGND VGND VPWR VPWR _12845_/Y sky130_fd_sc_hd__inv_2
X_15633_ _12585_/Y _15628_/X _15286_/X _15593_/A VGND VGND VPWR VPWR _24504_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18352_ _18352_/A VGND VGND VPWR VPWR _18491_/A sky130_fd_sc_hd__buf_2
X_12776_ _23013_/A VGND VGND VPWR VPWR _12890_/A sky130_fd_sc_hd__inv_2
X_15564_ _15562_/Y _15558_/X _15563_/X _15558_/X VGND VGND VPWR VPWR _15564_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20827__A _15637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _24393_/Q VGND VGND VPWR VPWR _17303_/Y sky130_fd_sc_hd__inv_2
XPHY_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11726_/Y VGND VGND VPWR VPWR _11960_/A sky130_fd_sc_hd__buf_2
X_14515_ _14501_/X _14505_/Y VGND VGND VPWR VPWR _14515_/Y sky130_fd_sc_hd__nor2_4
XPHY_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _15464_/X VGND VGND VPWR VPWR _15495_/X sky130_fd_sc_hd__buf_2
X_18283_ _18202_/Y _18277_/B VGND VGND VPWR VPWR _18283_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__14825__A _24155_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14843__A2_N _24144_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17234_ _17224_/Y _18095_/B _17226_/X _17233_/X VGND VGND VPWR VPWR _17234_/X sky130_fd_sc_hd__o22a_4
XPHY_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ _23925_/Q VGND VGND VPWR VPWR _22484_/A sky130_fd_sc_hd__inv_2
X_14446_ _14440_/X _14444_/B _14445_/Y VGND VGND VPWR VPWR _14446_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18016__B _13619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14377_ _14377_/A _14377_/B VGND VGND VPWR VPWR _14378_/A sky130_fd_sc_hd__and2_4
X_17165_ _17086_/X _17161_/X _17164_/Y VGND VGND VPWR VPWR _24029_/D sky130_fd_sc_hd__and3_4
XFILLER_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11589_ HWDATA[13] VGND VGND VPWR VPWR _16093_/A sky130_fd_sc_hd__buf_2
XANTENNA__23946__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13328_ _13328_/A VGND VGND VPWR VPWR _13328_/X sky130_fd_sc_hd__buf_2
X_16116_ _24328_/Q VGND VGND VPWR VPWR _16116_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14858__A2_N _14859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17096_ _17042_/X _17096_/B VGND VGND VPWR VPWR _17097_/B sky130_fd_sc_hd__or2_4
XFILLER_115_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15656__A _22147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13259_ _13120_/X _13259_/B VGND VGND VPWR VPWR _13259_/X sky130_fd_sc_hd__or2_4
X_16047_ _16037_/Y _16046_/X _15828_/X _16046_/X VGND VGND VPWR VPWR _24355_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12999__B _13008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19806_ _19800_/X _18067_/X _15704_/X _13170_/B _19802_/X VGND VGND VPWR VPWR _23203_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_9_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17998_ _17982_/X _17990_/X _15704_/X _23914_/Q _17983_/X VGND VGND VPWR VPWR _23914_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21393__A _21393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19737_ _19737_/A VGND VGND VPWR VPWR _19737_/Y sky130_fd_sc_hd__inv_2
X_16949_ _16832_/Y _16953_/A VGND VGND VPWR VPWR _16949_/Y sky130_fd_sc_hd__nand2_4
XFILLER_49_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13664__B1 _13663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19668_ _19680_/A VGND VGND VPWR VPWR _19668_/X sky130_fd_sc_hd__buf_2
XANTENNA__24734__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_8_0_HCLK clkbuf_4_4_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18619_ _18619_/A _18619_/B VGND VGND VPWR VPWR _18619_/X sky130_fd_sc_hd__or2_4
XANTENNA__22901__A1_N _12417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19599_ _19599_/A VGND VGND VPWR VPWR _21913_/B sky130_fd_sc_hd__inv_2
X_21630_ _21626_/A _21630_/B _21629_/X VGND VGND VPWR VPWR _21630_/X sky130_fd_sc_hd__and3_4
XANTENNA__16934__B _16927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21561_ _22279_/A VGND VGND VPWR VPWR _21561_/X sky130_fd_sc_hd__buf_2
X_23300_ _23939_/CLK _19540_/X VGND VGND VPWR VPWR _23300_/Q sky130_fd_sc_hd__dfxtp_4
X_20512_ _20512_/A VGND VGND VPWR VPWR _20512_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24280_ _24138_/CLK _16250_/X HRESETn VGND VGND VPWR VPWR _24280_/Q sky130_fd_sc_hd__dfrtp_4
X_21492_ _23105_/Q _21638_/A _23081_/Q _15642_/X VGND VGND VPWR VPWR _21492_/X sky130_fd_sc_hd__o22a_4
XFILLER_18_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23231_ _23383_/CLK _23231_/D VGND VGND VPWR VPWR _19733_/A sky130_fd_sc_hd__dfxtp_4
X_20443_ _21887_/A _13505_/B _20442_/Y VGND VGND VPWR VPWR _20443_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__22454__A2 _22451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19855__B1 _19832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23687__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16669__B1 _24097_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23162_ _23308_/CLK _19916_/X VGND VGND VPWR VPWR _19915_/A sky130_fd_sc_hd__dfxtp_4
X_20374_ _20374_/A _20372_/Y _20373_/X VGND VGND VPWR VPWR _20374_/X sky130_fd_sc_hd__and3_4
XANTENNA__23616__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22113_ _21339_/A _22105_/X _22112_/X VGND VGND VPWR VPWR _22113_/X sky130_fd_sc_hd__and3_4
XANTENNA__14144__A1 _20889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15566__A _15561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15341__B1 _11548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23093_ _23100_/CLK _20099_/X VGND VGND VPWR VPWR _23093_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_133_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22044_ _22041_/Y _22042_/X _22043_/X _23917_/Q _21400_/A VGND VGND VPWR VPWR _22044_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18877__A _18876_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22399__A _22399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_253_0_HCLK clkbuf_8_253_0_HCLK/A VGND VGND VPWR VPWR _24676_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_87_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23995_ _25214_/CLK _17390_/X HRESETn VGND VGND VPWR VPWR _17270_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21717__B2 _13618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22946_ _21175_/X _22944_/X _13362_/A _22945_/X VGND VGND VPWR VPWR _22946_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24475__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24404__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22877_ _14901_/A _22616_/X _22351_/X VGND VGND VPWR VPWR _22877_/X sky130_fd_sc_hd__o21a_4
X_12630_ _12739_/A _24508_/Q _12629_/X _24505_/Q VGND VGND VPWR VPWR _12630_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21828_ _20980_/A _21826_/X _21827_/X VGND VGND VPWR VPWR _21828_/X sky130_fd_sc_hd__and3_4
XANTENNA__21750__B _21251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24616_ _24587_/CLK _24616_/D HRESETn VGND VGND VPWR VPWR _24616_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14080__B1 _13663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22142__A1 _21707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20647__A _20647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11969__B1 _11616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _25058_/Q _12559_/Y _12547_/A _12560_/Y VGND VGND VPWR VPWR _12561_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23023__A _23023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24547_ _24521_/CLK _15524_/X HRESETn VGND VGND VPWR VPWR _24547_/Q sky130_fd_sc_hd__dfrtp_4
X_21759_ _21010_/A VGND VGND VPWR VPWR _21764_/A sky130_fd_sc_hd__buf_2
XANTENNA__20153__B1 _15416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12630__B2 _24505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11512_ _23759_/Q VGND VGND VPWR VPWR _11512_/Y sky130_fd_sc_hd__inv_2
X_14300_ _14288_/A VGND VGND VPWR VPWR _14300_/X sky130_fd_sc_hd__buf_2
XANTENNA__17021__A _17021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15280_ _15278_/Y _15276_/X _15279_/X _15276_/X VGND VGND VPWR VPWR _15280_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12492_ _12492_/A VGND VGND VPWR VPWR _25084_/D sky130_fd_sc_hd__inv_2
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24478_ _24478_/CLK _15694_/X HRESETn VGND VGND VPWR VPWR _24478_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14231_ HWDATA[6] VGND VGND VPWR VPWR _16373_/A sky130_fd_sc_hd__buf_2
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17248__A1_N _25211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23429_ _25067_/CLK _19173_/X VGND VGND VPWR VPWR _23429_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_138_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14162_ _24835_/Q _14161_/Y _12053_/A VGND VGND VPWR VPWR _14162_/X sky130_fd_sc_hd__o21a_4
XFILLER_137_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13113_ _13113_/A _13101_/X _13113_/C VGND VGND VPWR VPWR _13113_/X sky130_fd_sc_hd__and3_4
X_14093_ _24856_/Q VGND VGND VPWR VPWR _14093_/Y sky130_fd_sc_hd__inv_2
X_18970_ _18982_/A VGND VGND VPWR VPWR _18970_/X sky130_fd_sc_hd__buf_2
XFILLER_124_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_63_0_HCLK clkbuf_6_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_63_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_13044_ _13040_/X _13043_/X _13026_/X VGND VGND VPWR VPWR _13044_/X sky130_fd_sc_hd__o21a_4
X_17921_ _17889_/A _17921_/B _17920_/X VGND VGND VPWR VPWR _17922_/C sky130_fd_sc_hd__and3_4
XFILLER_3_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15195__B _15159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17852_ _17816_/A _23434_/Q VGND VGND VPWR VPWR _17852_/X sky130_fd_sc_hd__or2_4
X_16803_ _24417_/Q _16802_/Y _15857_/Y _24079_/Q VGND VGND VPWR VPWR _16803_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17783_ _17783_/A _17783_/B _17783_/C VGND VGND VPWR VPWR _17783_/X sky130_fd_sc_hd__and3_4
XANTENNA__13646__B1 _13645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14995_ _14995_/A _15094_/A VGND VGND VPWR VPWR _14995_/X sky130_fd_sc_hd__or2_4
XFILLER_47_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22102__A _20972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21708__A1 _18117_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21708__B2 _20747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19522_ _23305_/Q VGND VGND VPWR VPWR _19522_/Y sky130_fd_sc_hd__inv_2
X_16734_ _15991_/Y _23946_/Q _22910_/A _16733_/Y VGND VGND VPWR VPWR _16739_/B sky130_fd_sc_hd__a2bb2o_4
X_13946_ _13939_/Y _13945_/Y _13933_/A VGND VGND VPWR VPWR _13946_/X sky130_fd_sc_hd__and3_4
XFILLER_130_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16100__A _16100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19453_ _21657_/B _19449_/X _19452_/X _19449_/X VGND VGND VPWR VPWR _23331_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15399__B1 _15282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16665_ _14732_/Y _16663_/X _16369_/X _16663_/X VGND VGND VPWR VPWR _24100_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24145__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13877_ _14352_/A _14357_/B _13877_/C _13877_/D VGND VGND VPWR VPWR _13878_/D sky130_fd_sc_hd__or4_4
XFILLER_34_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18404_ _24218_/Q _18452_/C _16464_/Y _18419_/A VGND VGND VPWR VPWR _18404_/X sky130_fd_sc_hd__a2bb2o_4
X_15616_ _15611_/X _15599_/X _15501_/X _24515_/Q _15612_/X VGND VGND VPWR VPWR _24515_/D
+ sky130_fd_sc_hd__a32o_4
X_12828_ _25006_/Q _12826_/Y _25010_/Q _12827_/Y VGND VGND VPWR VPWR _12828_/X sky130_fd_sc_hd__a2bb2o_4
X_19384_ _19383_/Y _19378_/X _19360_/X _19378_/X VGND VGND VPWR VPWR _19384_/X sky130_fd_sc_hd__a2bb2o_4
X_16596_ _16594_/Y _16595_/X _15497_/X _16595_/X VGND VGND VPWR VPWR _16596_/X sky130_fd_sc_hd__a2bb2o_4
X_18335_ _18327_/B _18335_/B _18319_/X VGND VGND VPWR VPWR _18335_/X sky130_fd_sc_hd__and3_4
XFILLER_91_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15547_ _15544_/Y _15537_/X _15545_/X _15546_/X VGND VGND VPWR VPWR _24539_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20144__B1 _15520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12759_ _12739_/B _12759_/B _12755_/X VGND VGND VPWR VPWR _12759_/X sky130_fd_sc_hd__and3_4
XPHY_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24632__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18266_ _18268_/B VGND VGND VPWR VPWR _18266_/Y sky130_fd_sc_hd__inv_2
X_15478_ _15368_/X _15461_/X _15477_/X _24571_/Q _15466_/X VGND VGND VPWR VPWR _24571_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_30_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17217_ _24012_/Q VGND VGND VPWR VPWR _17217_/Y sky130_fd_sc_hd__inv_2
X_14429_ _11505_/A _20842_/B _11726_/Y _13609_/X VGND VGND VPWR VPWR _14429_/X sky130_fd_sc_hd__or4_4
X_18197_ _23875_/Q VGND VGND VPWR VPWR _18223_/A sky130_fd_sc_hd__inv_2
XANTENNA__12075__A _12075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17148_ _17145_/A _17145_/B VGND VGND VPWR VPWR _17148_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15386__A _16369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17079_ _17079_/A VGND VGND VPWR VPWR _17079_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20090_ _21332_/B _20089_/X _19614_/A _20089_/X VGND VGND VPWR VPWR _23096_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24986__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24915__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22800_ _22495_/A _22787_/Y _22800_/C _22799_/Y VGND VGND VPWR VPWR _22801_/D sky130_fd_sc_hd__or4_4
Xclkbuf_8_20_0_HCLK clkbuf_8_21_0_HCLK/A VGND VGND VPWR VPWR _24953_/CLK sky130_fd_sc_hd__clkbuf_1
X_23780_ _23100_/CLK _20685_/X HRESETn VGND VGND VPWR VPWR RsTx_S0 sky130_fd_sc_hd__dfstp_4
X_20992_ _21012_/A VGND VGND VPWR VPWR _20998_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_83_0_HCLK clkbuf_8_83_0_HCLK/A VGND VGND VPWR VPWR _24783_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_93_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21851__A _21851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22731_ _24049_/Q _22952_/B VGND VGND VPWR VPWR _22734_/B sky130_fd_sc_hd__or2_4
XFILLER_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20922__A2 _11940_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22662_ _11562_/Y _22536_/X _15950_/Y _22537_/X VGND VGND VPWR VPWR _22662_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22124__A1 _21178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22124__B2 _16393_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24401_ _24399_/CLK _15895_/X HRESETn VGND VGND VPWR VPWR _15892_/A sky130_fd_sc_hd__dfrtp_4
X_21613_ _21625_/A _19675_/Y VGND VGND VPWR VPWR _21613_/X sky130_fd_sc_hd__or2_4
XFILLER_80_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22855__A1_N _12416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22593_ _22702_/A _22592_/X VGND VGND VPWR VPWR _22593_/X sky130_fd_sc_hd__and2_4
XANTENNA__23868__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24332_ _23852_/CLK _24332_/D HRESETn VGND VGND VPWR VPWR _24332_/Q sky130_fd_sc_hd__dfrtp_4
X_21544_ _21544_/A VGND VGND VPWR VPWR _21544_/X sky130_fd_sc_hd__buf_2
XANTENNA__21883__B1 _24099_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17776__A _17716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24263_ _24662_/CLK _16283_/X HRESETn VGND VGND VPWR VPWR _24263_/Q sky130_fd_sc_hd__dfrtp_4
X_21475_ _21342_/A _21475_/B VGND VGND VPWR VPWR _21475_/X sky130_fd_sc_hd__or2_4
X_23214_ _23308_/CLK _23214_/D VGND VGND VPWR VPWR _23214_/Q sky130_fd_sc_hd__dfxtp_4
X_20426_ _13498_/Y _13499_/Y _13501_/Y VGND VGND VPWR VPWR _20426_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21298__A _14747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24194_ _24225_/CLK _24194_/D HRESETn VGND VGND VPWR VPWR _24194_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15296__A HTRANS[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23145_ _25044_/CLK _19961_/X VGND VGND VPWR VPWR _23145_/Q sky130_fd_sc_hd__dfxtp_4
X_20357_ _14618_/A VGND VGND VPWR VPWR _20357_/X sky130_fd_sc_hd__buf_2
XFILLER_49_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16657__A3 _16096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23076_ _23993_/CLK _23076_/D VGND VGND VPWR VPWR _23076_/Q sky130_fd_sc_hd__dfxtp_4
X_20288_ _20288_/A _20283_/A VGND VGND VPWR VPWR _20288_/Y sky130_fd_sc_hd__nand2_4
X_22027_ _13934_/A _21544_/A _23617_/Q _22218_/C VGND VGND VPWR VPWR _22027_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24656__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13800_ _13800_/A _13800_/B VGND VGND VPWR VPWR _13800_/X sky130_fd_sc_hd__or2_4
XFILLER_91_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14245__A1_N _14004_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11992_ _11992_/A VGND VGND VPWR VPWR _11992_/Y sky130_fd_sc_hd__inv_2
X_14780_ _14880_/A _22857_/A _24702_/Q _14779_/Y VGND VGND VPWR VPWR _14784_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23978_ _23979_/CLK _23978_/D HRESETn VGND VGND VPWR VPWR _23978_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_44_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22857__A _22857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13731_ _24637_/Q VGND VGND VPWR VPWR _13732_/D sky130_fd_sc_hd__inv_2
X_22929_ _16054_/A _22311_/A _22864_/X VGND VGND VPWR VPWR _22929_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16855__A _16774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20913__A2 _14016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16450_ _16450_/A VGND VGND VPWR VPWR _16450_/Y sky130_fd_sc_hd__inv_2
X_13662_ _13437_/Y _13657_/X _11607_/X _13661_/X VGND VGND VPWR VPWR _13662_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15401_ _15401_/A VGND VGND VPWR VPWR _15401_/X sky130_fd_sc_hd__buf_2
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12613_ _12612_/Y _12619_/A _12648_/A _12556_/Y VGND VGND VPWR VPWR _12613_/X sky130_fd_sc_hd__a2bb2o_4
X_13593_ _13559_/A _13559_/B VGND VGND VPWR VPWR _13593_/Y sky130_fd_sc_hd__nand2_4
X_16381_ _16381_/A VGND VGND VPWR VPWR _16381_/Y sky130_fd_sc_hd__inv_2
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18120_ _18120_/A VGND VGND VPWR VPWR _21586_/B sky130_fd_sc_hd__inv_2
XFILLER_101_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12544_ _25068_/Q VGND VGND VPWR VPWR _12544_/Y sky130_fd_sc_hd__inv_2
X_15332_ HWDATA[28] VGND VGND VPWR VPWR _15332_/X sky130_fd_sc_hd__buf_2
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18051_ _23903_/Q VGND VGND VPWR VPWR _20034_/A sky130_fd_sc_hd__buf_2
X_12475_ _12412_/C _12480_/B _12427_/X VGND VGND VPWR VPWR _12475_/Y sky130_fd_sc_hd__a21oi_4
X_15263_ _13730_/X _15260_/X _15256_/X _13728_/X _15262_/X VGND VGND VPWR VPWR _15263_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16590__A _16566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17002_ _16174_/Y _16992_/A _24310_/Q _16968_/Y VGND VGND VPWR VPWR _17004_/C sky130_fd_sc_hd__a2bb2o_4
X_14214_ _14211_/Y _14212_/X _14213_/X _14202_/X VGND VGND VPWR VPWR _14214_/X sky130_fd_sc_hd__a2bb2o_4
X_15194_ _15193_/X VGND VGND VPWR VPWR _24662_/D sky130_fd_sc_hd__inv_2
XFILLER_67_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14145_ _12053_/Y VGND VGND VPWR VPWR _14145_/X sky130_fd_sc_hd__buf_2
XANTENNA__16648__A3 HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15305__B1 HADDR[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14076_ _14070_/Y _14075_/Y sda_oen_o_S5 _14070_/Y VGND VGND VPWR VPWR _14076_/X
+ sky130_fd_sc_hd__a2bb2o_4
X_18953_ _16545_/X VGND VGND VPWR VPWR _18953_/X sky130_fd_sc_hd__buf_2
XFILLER_80_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19751__A2_N _19750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13027_ _13018_/X _13024_/X _13026_/X VGND VGND VPWR VPWR _13027_/X sky130_fd_sc_hd__o21a_4
X_17904_ _17968_/A _17904_/B _17903_/X VGND VGND VPWR VPWR _17904_/X sky130_fd_sc_hd__and3_4
X_18884_ _18876_/Y VGND VGND VPWR VPWR _18884_/X sky130_fd_sc_hd__buf_2
XANTENNA__24397__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16805__B1 _24396_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17835_ _17961_/A _17833_/X _17834_/X VGND VGND VPWR VPWR _17835_/X sky130_fd_sc_hd__and3_4
XFILLER_39_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24326__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17766_ _15730_/X _17739_/X _17764_/X _23933_/Q _17765_/X VGND VGND VPWR VPWR _17766_/X
+ sky130_fd_sc_hd__o32a_4
X_14978_ _14980_/B VGND VGND VPWR VPWR _14979_/B sky130_fd_sc_hd__inv_2
X_19505_ _23311_/Q VGND VGND VPWR VPWR _19505_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16717_ _16717_/A _16717_/B _16707_/X _16716_/X VGND VGND VPWR VPWR _16746_/A sky130_fd_sc_hd__or4_4
X_13929_ _24890_/Q _13928_/X _24891_/Q VGND VGND VPWR VPWR _13930_/B sky130_fd_sc_hd__or3_4
X_17697_ _17697_/A _17697_/B VGND VGND VPWR VPWR _17697_/X sky130_fd_sc_hd__or2_4
XFILLER_63_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20904__A2 _20826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22486__B _22486_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19436_ _23335_/Q VGND VGND VPWR VPWR _19436_/Y sky130_fd_sc_hd__inv_2
X_16648_ _16624_/X _16625_/X HWDATA[16] _22502_/A _16647_/X VGND VGND VPWR VPWR _16648_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14044__B1 _13635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19367_ _19365_/Y _19363_/X _19366_/X _19363_/X VGND VGND VPWR VPWR _23360_/D sky130_fd_sc_hd__a2bb2o_4
X_16579_ _15799_/X _16573_/X _15596_/X _24150_/Q _16566_/X VGND VGND VPWR VPWR _24150_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_22_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15792__B1 _15513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23961__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18318_ _18318_/A _18302_/X VGND VGND VPWR VPWR _18320_/B sky130_fd_sc_hd__nand2_4
XANTENNA__25185__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19298_ _19298_/A VGND VGND VPWR VPWR _19298_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25114__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18249_ _18249_/A VGND VGND VPWR VPWR _18249_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19704__A2_N _19701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21260_ _13630_/C VGND VGND VPWR VPWR _21793_/A sky130_fd_sc_hd__buf_2
X_20211_ _20204_/X VGND VGND VPWR VPWR _20212_/B sky130_fd_sc_hd__buf_2
XANTENNA__13629__A _16042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21191_ _11720_/X VGND VGND VPWR VPWR _22045_/B sky130_fd_sc_hd__inv_2
XFILLER_116_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20840__A1 _12793_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20142_ _20140_/Y _20136_/X _13668_/A _20141_/X VGND VGND VPWR VPWR _23074_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19719__A2_N _19710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20750__A _20749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15844__A _24420_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20073_ _20072_/Y _20067_/X _15416_/X _20067_/X VGND VGND VPWR VPWR _20073_/X sky130_fd_sc_hd__a2bb2o_4
X_24950_ _24957_/CLK _24950_/D HRESETn VGND VGND VPWR VPWR _11663_/A sky130_fd_sc_hd__dfrtp_4
X_23901_ _23343_/CLK _18040_/X HRESETn VGND VGND VPWR VPWR _23901_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24067__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24881_ _23648_/CLK _24881_/D HRESETn VGND VGND VPWR VPWR _13925_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_22_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23832_ _23830_/CLK _23832_/D HRESETn VGND VGND VPWR VPWR _23832_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14283__B1 _14094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22677__A _22677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21581__A _21581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23763_ _24013_/CLK _20197_/X HRESETn VGND VGND VPWR VPWR _23763_/Q sky130_fd_sc_hd__dfrtp_4
X_20975_ _20975_/A _20975_/B _20974_/X VGND VGND VPWR VPWR _20975_/X sky130_fd_sc_hd__and3_4
XFILLER_72_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22714_ _16692_/A _22654_/X _22608_/X VGND VGND VPWR VPWR _22716_/C sky130_fd_sc_hd__a21o_4
XANTENNA__14035__B1 _13632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23694_ _23668_/CLK _20238_/X HRESETn VGND VGND VPWR VPWR _23694_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20108__B1 _19610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22645_ _24308_/Q _22897_/B VGND VGND VPWR VPWR _22645_/X sky130_fd_sc_hd__or2_4
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11612__A _13663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22576_ _22576_/A VGND VGND VPWR VPWR _22576_/X sky130_fd_sc_hd__buf_2
XFILLER_51_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23631__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21320__A2 _15456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21527_ _21523_/X _21526_/X _21242_/X VGND VGND VPWR VPWR _21528_/C sky130_fd_sc_hd__o21a_4
XFILLER_103_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24315_ _24049_/CLK _24315_/D HRESETn VGND VGND VPWR VPWR _24315_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12260_ _12132_/Y _12257_/X VGND VGND VPWR VPWR _12260_/X sky130_fd_sc_hd__or2_4
X_24246_ _24213_/CLK _16327_/X HRESETn VGND VGND VPWR VPWR _16325_/A sky130_fd_sc_hd__dfrtp_4
X_21458_ _21458_/A _21428_/Y _21434_/X _21457_/X VGND VGND VPWR VPWR _21458_/X sky130_fd_sc_hd__or4_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23020__B _23020_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15738__B _15741_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20409_ _13800_/A _20205_/Y _20409_/C VGND VGND VPWR VPWR _20410_/A sky130_fd_sc_hd__or3_4
X_12191_ _12186_/B _12423_/A VGND VGND VPWR VPWR _12192_/B sky130_fd_sc_hd__and2_4
X_24177_ _24177_/CLK _16509_/X HRESETn VGND VGND VPWR VPWR _24177_/Q sky130_fd_sc_hd__dfrtp_4
X_21389_ _21227_/A _21389_/B VGND VGND VPWR VPWR _21391_/B sky130_fd_sc_hd__or2_4
XFILLER_123_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23128_ _23128_/CLK _23128_/D VGND VGND VPWR VPWR _13262_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_134_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15950_ _24380_/Q VGND VGND VPWR VPWR _15950_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23059_ _20737_/X VGND VGND VPWR VPWR IRQ[7] sky130_fd_sc_hd__buf_2
XANTENNA__24490__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18788__B1 _18740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14901_ _14901_/A VGND VGND VPWR VPWR _14901_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15881_ _15879_/Y _15880_/X _11598_/X _15880_/X VGND VGND VPWR VPWR _24406_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17620_ _17614_/A _17614_/B VGND VGND VPWR VPWR _17620_/Y sky130_fd_sc_hd__nand2_4
XFILLER_48_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14832_ _24687_/Q _14801_/Y _24692_/Q _14831_/Y VGND VGND VPWR VPWR _14832_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14274__B1 _14236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21491__A _21491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17551_ _17497_/D _17550_/X VGND VGND VPWR VPWR _17554_/B sky130_fd_sc_hd__or2_4
X_14763_ _14762_/Y VGND VGND VPWR VPWR _15019_/A sky130_fd_sc_hd__buf_2
X_11975_ _11975_/A VGND VGND VPWR VPWR _11975_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16502_ _16501_/Y _16499_/X _16254_/X _16499_/X VGND VGND VPWR VPWR _24180_/D sky130_fd_sc_hd__a2bb2o_4
X_13714_ _13754_/B VGND VGND VPWR VPWR _13742_/C sky130_fd_sc_hd__buf_2
XFILLER_17_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17482_ _17482_/A VGND VGND VPWR VPWR _17483_/A sky130_fd_sc_hd__inv_2
X_14694_ _14694_/A VGND VGND VPWR VPWR _14869_/A sky130_fd_sc_hd__inv_2
XANTENNA__23719__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19221_ _11625_/A VGND VGND VPWR VPWR _19221_/X sky130_fd_sc_hd__buf_2
XANTENNA__18960__B1 _18959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16433_ _16401_/A VGND VGND VPWR VPWR _16452_/A sky130_fd_sc_hd__buf_2
X_13645_ _14218_/A VGND VGND VPWR VPWR _13645_/X sky130_fd_sc_hd__buf_2
XANTENNA__15774__B1 _15772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11522__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19152_ _18743_/X VGND VGND VPWR VPWR _19152_/X sky130_fd_sc_hd__buf_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16364_ _16364_/A VGND VGND VPWR VPWR _16364_/X sky130_fd_sc_hd__buf_2
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ _13550_/Y VGND VGND VPWR VPWR _13576_/X sky130_fd_sc_hd__buf_2
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ _18099_/Y _18102_/Y _18099_/A _18101_/X VGND VGND VPWR VPWR _23889_/D sky130_fd_sc_hd__o22a_4
X_15315_ _11949_/A _14195_/B _14195_/C _15314_/X VGND VGND VPWR VPWR _15315_/X sky130_fd_sc_hd__or4_4
XANTENNA__21311__A1_N _14259_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12527_ _12379_/Y _12502_/X _12444_/A _12525_/B VGND VGND VPWR VPWR _12527_/X sky130_fd_sc_hd__a211o_4
X_19083_ _23460_/Q VGND VGND VPWR VPWR _19083_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15526__B1 _24545_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16295_ _16294_/Y _16247_/A _16219_/X _16247_/A VGND VGND VPWR VPWR _24255_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20554__B _20554_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18034_ _18023_/A _18033_/X VGND VGND VPWR VPWR _18034_/X sky130_fd_sc_hd__and2_4
X_15246_ _13776_/C _14100_/X _15240_/X _13753_/A _15245_/X VGND VGND VPWR VPWR _24648_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_8_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13001__A1 _12858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12458_ _12458_/A VGND VGND VPWR VPWR _12458_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15648__B _15459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19807__A3 _18000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21075__B2 _22018_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12389_ _12388_/Y VGND VGND VPWR VPWR _12389_/X sky130_fd_sc_hd__buf_2
X_15177_ _15177_/A _15177_/B VGND VGND VPWR VPWR _15177_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24578__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14128_ MSO_S2 _14127_/X _24847_/Q _14122_/X VGND VGND VPWR VPWR _14128_/Y sky130_fd_sc_hd__a22oi_4
X_19985_ _21233_/B _19982_/X _15561_/X _19982_/X VGND VGND VPWR VPWR _19985_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24507__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15664__A _15664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14059_ _14059_/A VGND VGND VPWR VPWR _14059_/Y sky130_fd_sc_hd__inv_2
X_18936_ _18934_/Y _18935_/X _18823_/X _18935_/X VGND VGND VPWR VPWR _23513_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14501__B2 _14484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18779__B1 _18685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18867_ _18865_/Y _18866_/X _18823_/X _18866_/X VGND VGND VPWR VPWR _18867_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24160__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18975__A _18982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13184__A _13102_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17818_ _17780_/A _17818_/B _17818_/C VGND VGND VPWR VPWR _17823_/B sky130_fd_sc_hd__and3_4
X_18798_ _18798_/A VGND VGND VPWR VPWR _18798_/X sky130_fd_sc_hd__buf_2
XANTENNA__14265__B1 _14218_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22497__A _16515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22327__B2 _20926_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17749_ _14577_/X VGND VGND VPWR VPWR _17935_/A sky130_fd_sc_hd__buf_2
XANTENNA__17203__B1 _17202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20760_ _20759_/X VGND VGND VPWR VPWR _21357_/A sky130_fd_sc_hd__buf_2
XFILLER_39_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19419_ _19415_/Y _19418_/X _19329_/X _19418_/X VGND VGND VPWR VPWR _19419_/X sky130_fd_sc_hd__a2bb2o_4
X_20691_ _20691_/A _20691_/B VGND VGND VPWR VPWR _23788_/D sky130_fd_sc_hd__and2_4
Xclkbuf_8_157_0_HCLK clkbuf_7_78_0_HCLK/X VGND VGND VPWR VPWR _24502_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22430_ _15655_/A VGND VGND VPWR VPWR _22505_/A sky130_fd_sc_hd__buf_2
XFILLER_91_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20745__A _20744_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15780__A3 _15494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18703__B1 _18679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22361_ _15970_/A _21543_/A VGND VGND VPWR VPWR _22361_/X sky130_fd_sc_hd__or2_4
XANTENNA__15517__B1 _15390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15839__A _24422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21853__A3 _22629_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23665__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24100_ _24101_/CLK _24100_/D HRESETn VGND VGND VPWR VPWR _14732_/A sky130_fd_sc_hd__dfrtp_4
X_21312_ _24794_/Q _20931_/X _21309_/X _21310_/X _21311_/X VGND VGND VPWR VPWR _21312_/X
+ sky130_fd_sc_hd__a2111o_4
X_25080_ _25097_/CLK _25080_/D HRESETn VGND VGND VPWR VPWR _25080_/Q sky130_fd_sc_hd__dfrtp_4
X_22292_ _22274_/Y _22495_/A _22292_/C _22292_/D VGND VGND VPWR VPWR _22292_/X sky130_fd_sc_hd__or4_4
XFILLER_15_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15532__A3 _15432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24031_ _24031_/CLK _24031_/D HRESETn VGND VGND VPWR VPWR _17027_/A sky130_fd_sc_hd__dfrtp_4
X_21243_ _21236_/X _21241_/X _21242_/X VGND VGND VPWR VPWR _21243_/X sky130_fd_sc_hd__o21a_4
XANTENNA__11686__A2_N _22215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24930__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21174_ _17636_/X _21162_/X _21174_/C VGND VGND VPWR VPWR _21174_/X sky130_fd_sc_hd__or3_4
XANTENNA__24248__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20125_ _17982_/A _20119_/X _18000_/X _23081_/Q _20117_/X VGND VGND VPWR VPWR _20125_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_132_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_22_0_HCLK_A clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15574__A _16624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22566__A1 _24562_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20056_ _20054_/X _15410_/X _13663_/A _22043_/A _20055_/X VGND VGND VPWR VPWR _20056_/X
+ sky130_fd_sc_hd__a32o_4
X_24933_ _24974_/CLK _13662_/X HRESETn VGND VGND VPWR VPWR _24933_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20577__B1 _20562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11607__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24864_ _24870_/CLK _14065_/X HRESETn VGND VGND VPWR VPWR _14064_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__14256__B1 _14209_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23815_ _23824_/CLK _23815_/D HRESETn VGND VGND VPWR VPWR _23815_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24795_ _24859_/CLK _24795_/D HRESETn VGND VGND VPWR VPWR _24795_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23883__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11759_/X VGND VGND VPWR VPWR _11760_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_53_0_HCLK clkbuf_6_26_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_53_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20958_ _20964_/A _20093_/Y VGND VGND VPWR VPWR _20958_/X sky130_fd_sc_hd__or2_4
XPHY_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23746_ _24177_/CLK _20642_/Y HRESETn VGND VGND VPWR VPWR _23746_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23812__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25036__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _23923_/Q VGND VGND VPWR VPWR _11691_/Y sky130_fd_sc_hd__inv_2
XPHY_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ _20889_/A _20759_/X VGND VGND VPWR VPWR _20889_/X sky130_fd_sc_hd__and2_4
XANTENNA__21740__A2_N _20818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23677_ _24728_/CLK _20392_/Y HRESETn VGND VGND VPWR VPWR _20389_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13430_ _13428_/A _14414_/A _13428_/Y _13429_/Y VGND VGND VPWR VPWR _13430_/X sky130_fd_sc_hd__o22a_4
XFILLER_41_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21829__B1 _21172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22628_ _24486_/Q _22757_/B VGND VGND VPWR VPWR _22628_/X sky130_fd_sc_hd__or2_4
XFILLER_42_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ _22745_/B VGND VGND VPWR VPWR _13362_/A sky130_fd_sc_hd__buf_2
XANTENNA__15508__B1 _24556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22559_ _15653_/X VGND VGND VPWR VPWR _22957_/B sky130_fd_sc_hd__buf_2
XFILLER_127_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15100_ _15159_/A VGND VGND VPWR VPWR _15123_/A sky130_fd_sc_hd__buf_2
X_12312_ _12312_/A _12312_/B _12312_/C _12312_/D VGND VGND VPWR VPWR _12312_/X sky130_fd_sc_hd__or4_4
X_13292_ _11751_/X _13290_/X _13292_/C VGND VGND VPWR VPWR _13292_/X sky130_fd_sc_hd__and3_4
X_16080_ _16080_/A VGND VGND VPWR VPWR _16080_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15523__A3 _15522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12243_ _12174_/B _12243_/B VGND VGND VPWR VPWR _12244_/B sky130_fd_sc_hd__or2_4
X_15031_ _14736_/X _15036_/B _14984_/X VGND VGND VPWR VPWR _15031_/Y sky130_fd_sc_hd__a21oi_4
X_24229_ _24197_/CLK _24229_/D HRESETn VGND VGND VPWR VPWR _24229_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24671__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20804__A1 _22014_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12174_ _12174_/A _12174_/B _12173_/X VGND VGND VPWR VPWR _12175_/C sky130_fd_sc_hd__or3_4
XFILLER_68_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20804__B2 _21591_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24600__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15484__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19770_ _21463_/B _19765_/X _19724_/X _19765_/X VGND VGND VPWR VPWR _19770_/X sky130_fd_sc_hd__a2bb2o_4
X_16982_ _24046_/Q VGND VGND VPWR VPWR _16982_/Y sky130_fd_sc_hd__inv_2
X_18721_ _18721_/A VGND VGND VPWR VPWR _18721_/Y sky130_fd_sc_hd__inv_2
X_15933_ _24387_/Q VGND VGND VPWR VPWR _15933_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20568__B1 _20562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18795__A _18678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18652_ _23611_/Q VGND VGND VPWR VPWR _18652_/Y sky130_fd_sc_hd__inv_2
X_15864_ _24412_/Q VGND VGND VPWR VPWR _15864_/Y sky130_fd_sc_hd__inv_2
X_17603_ _17603_/A _17603_/B _17602_/Y VGND VGND VPWR VPWR _17603_/X sky130_fd_sc_hd__and3_4
X_14815_ _24711_/Q _14814_/A _14990_/A _14814_/Y VGND VGND VPWR VPWR _14820_/B sky130_fd_sc_hd__o22a_4
X_18583_ _16375_/A _18421_/B _24232_/Q _18425_/A VGND VGND VPWR VPWR _18583_/X sky130_fd_sc_hd__a2bb2o_4
X_15795_ _15767_/X VGND VGND VPWR VPWR _15795_/X sky130_fd_sc_hd__buf_2
XFILLER_40_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22110__A _20966_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17534_ _16702_/Y _17534_/B VGND VGND VPWR VPWR _17535_/A sky130_fd_sc_hd__or2_4
X_14746_ _24684_/Q VGND VGND VPWR VPWR _15087_/A sky130_fd_sc_hd__inv_2
X_11958_ _11936_/Y _11957_/Y _11643_/X _11957_/Y VGND VGND VPWR VPWR _11958_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18933__B1 _18932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17465_ _17465_/A VGND VGND VPWR VPWR _17465_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15747__B1 _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14677_ _14633_/X _14610_/B _24718_/Q _14676_/X VGND VGND VPWR VPWR _14677_/X sky130_fd_sc_hd__a2bb2o_4
X_11889_ _11881_/A _11881_/B _11888_/Y VGND VGND VPWR VPWR _11891_/A sky130_fd_sc_hd__o21a_4
X_19204_ _19196_/A VGND VGND VPWR VPWR _19204_/X sky130_fd_sc_hd__buf_2
X_16416_ _24213_/Q VGND VGND VPWR VPWR _16416_/Y sky130_fd_sc_hd__inv_2
X_13628_ _22018_/B VGND VGND VPWR VPWR _16042_/A sky130_fd_sc_hd__buf_2
X_17396_ _17311_/Y _17371_/X _17345_/X _17393_/Y VGND VGND VPWR VPWR _17396_/X sky130_fd_sc_hd__a211o_4
XFILLER_34_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12067__B _16302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19135_ _19134_/Y _19130_/X _19089_/X _19130_/X VGND VGND VPWR VPWR _19135_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16347_ _16364_/A VGND VGND VPWR VPWR _16347_/X sky130_fd_sc_hd__buf_2
XANTENNA__15659__A _16305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13559_ _13559_/A _13559_/B VGND VGND VPWR VPWR _13559_/X sky130_fd_sc_hd__or2_4
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24759__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12981__B1 _12922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19066_ _17812_/B VGND VGND VPWR VPWR _19066_/Y sky130_fd_sc_hd__inv_2
X_16278_ _16262_/A VGND VGND VPWR VPWR _16278_/X sky130_fd_sc_hd__buf_2
XFILLER_103_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18017_ _17999_/X _15657_/X _11643_/A _23904_/Q _18016_/X VGND VGND VPWR VPWR _23904_/D
+ sky130_fd_sc_hd__a32o_4
X_15229_ _15229_/A VGND VGND VPWR VPWR _15230_/B sky130_fd_sc_hd__inv_2
XFILLER_114_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22796__A1 _12101_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19110__B1 _19109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22796__B2 _22238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21396__A _21396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24341__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19968_ _14493_/X _19862_/B _19509_/C VGND VGND VPWR VPWR _19969_/A sky130_fd_sc_hd__or3_4
XFILLER_101_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13289__B2 _13054_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22004__B _21907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18919_ _17684_/B VGND VGND VPWR VPWR _18919_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19899_ _19899_/A VGND VGND VPWR VPWR _21221_/B sky130_fd_sc_hd__inv_2
XFILLER_132_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21930_ _21930_/A _21926_/X _21929_/X VGND VGND VPWR VPWR _21930_/X sky130_fd_sc_hd__or3_4
XFILLER_83_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14238__B1 _14236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21861_ _22226_/A _21860_/X _14836_/Y _20757_/X VGND VGND VPWR VPWR _21861_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14789__B2 _24097_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20812_ _22564_/B VGND VGND VPWR VPWR _22429_/B sky130_fd_sc_hd__buf_2
X_23600_ _23992_/CLK _23600_/D VGND VGND VPWR VPWR _18684_/A sky130_fd_sc_hd__dfxtp_4
X_21792_ _11964_/A _21749_/X _21758_/Y _21642_/X _21791_/X VGND VGND VPWR VPWR _21792_/X
+ sky130_fd_sc_hd__a32o_4
X_24580_ _25183_/CLK _24580_/D HRESETn VGND VGND VPWR VPWR _14434_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22955__A _22167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22720__B2 _22029_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20743_ _21113_/C VGND VGND VPWR VPWR _20800_/A sky130_fd_sc_hd__buf_2
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23531_ _23531_/CLK _23531_/D VGND VGND VPWR VPWR _23531_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23462_ _23457_/CLK _23462_/D VGND VGND VPWR VPWR _17677_/B sky130_fd_sc_hd__dfxtp_4
X_20674_ _20556_/X _20673_/Y _16485_/A _20602_/X VGND VGND VPWR VPWR _23755_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22413_ _16441_/Y _21882_/X _16655_/Y _22017_/X VGND VGND VPWR VPWR _22413_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21287__A1 _22610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25201_ _23969_/CLK _11600_/X HRESETn VGND VGND VPWR VPWR _25201_/Q sky130_fd_sc_hd__dfrtp_4
X_23393_ _23411_/CLK _23393_/D VGND VGND VPWR VPWR _23393_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22344_ _22344_/A _16393_/D VGND VGND VPWR VPWR _22344_/X sky130_fd_sc_hd__and2_4
X_25132_ _25084_/CLK _12197_/Y HRESETn VGND VGND VPWR VPWR _12154_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_128_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16163__B1 _15765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24429__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25063_ _25061_/CLK _12686_/Y HRESETn VGND VGND VPWR VPWR _25063_/Q sky130_fd_sc_hd__dfrtp_4
X_22275_ _21581_/A _21300_/B _11950_/X _22510_/B VGND VGND VPWR VPWR _22275_/X sky130_fd_sc_hd__or4_4
XANTENNA__12724__B1 _12674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24014_ _24013_/CLK _24014_/D HRESETn VGND VGND VPWR VPWR _24014_/Q sky130_fd_sc_hd__dfrtp_4
X_21226_ _14443_/B VGND VGND VPWR VPWR _21227_/A sky130_fd_sc_hd__buf_2
XANTENNA__24082__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21157_ _17629_/B VGND VGND VPWR VPWR _21158_/A sky130_fd_sc_hd__buf_2
XANTENNA__24011__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20108_ _21474_/B _20103_/X _19610_/A _20103_/X VGND VGND VPWR VPWR _23089_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21088_ _21088_/A VGND VGND VPWR VPWR _21088_/X sky130_fd_sc_hd__buf_2
XFILLER_8_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12930_ _12883_/X _12892_/X _12845_/Y VGND VGND VPWR VPWR _12930_/X sky130_fd_sc_hd__o21a_4
X_20039_ _21932_/B _20036_/X _19714_/X _20036_/X VGND VGND VPWR VPWR _23116_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24916_ _24923_/CLK _13705_/X HRESETn VGND VGND VPWR VPWR _24916_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14229__B1 _14228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13255__C _13254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19535__A2_N _19534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25217__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12861_ _12860_/Y _24459_/Q _12860_/Y _24459_/Q VGND VGND VPWR VPWR _12865_/B sky130_fd_sc_hd__a2bb2o_4
X_24847_ _24847_/CLK _24847_/D HRESETn VGND VGND VPWR VPWR _24847_/Q sky130_fd_sc_hd__dfrtp_4
X_14600_ _19123_/D _14598_/Y _19123_/B _16035_/B VGND VGND VPWR VPWR _24733_/D sky130_fd_sc_hd__o22a_4
X_11812_ _11782_/X _11802_/A _11811_/Y VGND VGND VPWR VPWR _11817_/B sky130_fd_sc_hd__o21a_4
X_15580_ _15741_/B VGND VGND VPWR VPWR _15740_/A sky130_fd_sc_hd__inv_2
X_12792_ _22712_/A _12790_/Y _22900_/A _12791_/Y VGND VGND VPWR VPWR _12795_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24778_ _23618_/CLK _14334_/X HRESETn VGND VGND VPWR VPWR _24778_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14367__B HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14531_ _21202_/A VGND VGND VPWR VPWR _21376_/A sky130_fd_sc_hd__buf_2
XPHY_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11743_/A VGND VGND VPWR VPWR _18085_/A sky130_fd_sc_hd__buf_2
XFILLER_14_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23729_ _24161_/CLK _23729_/D HRESETn VGND VGND VPWR VPWR _13525_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _17250_/A _17245_/X _17248_/X _17249_/X VGND VGND VPWR VPWR _17269_/B sky130_fd_sc_hd__or4_4
XPHY_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14524_/A _14461_/X _14524_/A _14461_/X VGND VGND VPWR VPWR _14462_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _23920_/Q VGND VGND VPWR VPWR _22272_/A sky130_fd_sc_hd__inv_2
XFILLER_53_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_140_0_HCLK clkbuf_7_70_0_HCLK/X VGND VGND VPWR VPWR _23425_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16201_ _16200_/Y _16196_/X _15890_/X _16196_/X VGND VGND VPWR VPWR _24296_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ _13413_/A VGND VGND VPWR VPWR _13413_/Y sky130_fd_sc_hd__inv_2
XPHY_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17181_ _20389_/A _20389_/B VGND VGND VPWR VPWR _17182_/B sky130_fd_sc_hd__or2_4
XANTENNA__22475__B1 _24042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15479__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14393_ _14392_/X VGND VGND VPWR VPWR _14393_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24852__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16132_ _15421_/X _16135_/B _15912_/X _24321_/Q _16131_/X VGND VGND VPWR VPWR _24321_/D
+ sky130_fd_sc_hd__a32o_4
X_13344_ _13338_/Y VGND VGND VPWR VPWR _13344_/X sky130_fd_sc_hd__buf_2
XANTENNA__16154__B1 _16153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16063_ _16063_/A VGND VGND VPWR VPWR _16063_/Y sky130_fd_sc_hd__inv_2
X_13275_ _13171_/A _13273_/X _13275_/C VGND VGND VPWR VPWR _13279_/B sky130_fd_sc_hd__and3_4
XANTENNA__15901__B1 _15279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14704__B2 _24118_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15014_ _15014_/A _15014_/B _15013_/X VGND VGND VPWR VPWR _24705_/D sky130_fd_sc_hd__and3_4
X_12226_ _12225_/X VGND VGND VPWR VPWR _25124_/D sky130_fd_sc_hd__inv_2
X_12157_ _25108_/Q VGND VGND VPWR VPWR _12157_/Y sky130_fd_sc_hd__inv_2
X_19822_ _19831_/A VGND VGND VPWR VPWR _19822_/X sky130_fd_sc_hd__buf_2
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12088_ _12088_/A VGND VGND VPWR VPWR _12088_/Y sky130_fd_sc_hd__inv_2
X_16965_ _16176_/Y _17041_/A _16176_/Y _17041_/A VGND VGND VPWR VPWR _16965_/X sky130_fd_sc_hd__a2bb2o_4
X_19753_ _21166_/B _19750_/X _19731_/X _19750_/X VGND VGND VPWR VPWR _19753_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15916_ _15916_/A _15422_/A VGND VGND VPWR VPWR _15916_/X sky130_fd_sc_hd__or2_4
X_18704_ _13234_/B VGND VGND VPWR VPWR _18704_/Y sky130_fd_sc_hd__inv_2
X_19684_ _19684_/A VGND VGND VPWR VPWR _19684_/Y sky130_fd_sc_hd__inv_2
X_16896_ _16765_/Y _16895_/X _16849_/X VGND VGND VPWR VPWR _16896_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__23734__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18635_ _11708_/A _11697_/Y _11696_/X VGND VGND VPWR VPWR _23803_/D sky130_fd_sc_hd__o21ai_4
X_15847_ _15847_/A VGND VGND VPWR VPWR _15847_/X sky130_fd_sc_hd__buf_2
XFILLER_64_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13462__A _13462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18566_ _18562_/X _18566_/B _18564_/X _18565_/X VGND VGND VPWR VPWR _18582_/A sky130_fd_sc_hd__or4_4
X_15778_ _12823_/Y _15773_/X _15777_/X _15773_/X VGND VGND VPWR VPWR _24446_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17517_ _16710_/A _17517_/B VGND VGND VPWR VPWR _17517_/X sky130_fd_sc_hd__or2_4
X_14729_ _24117_/Q VGND VGND VPWR VPWR _14729_/Y sky130_fd_sc_hd__inv_2
X_18497_ _18434_/C _18501_/B _18496_/Y VGND VGND VPWR VPWR _23832_/D sky130_fd_sc_hd__o21a_4
XFILLER_21_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17448_ _17448_/A _17448_/B _21363_/A _11828_/X VGND VGND VPWR VPWR _17460_/B sky130_fd_sc_hd__or4_4
XFILLER_33_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17379_ _17378_/X VGND VGND VPWR VPWR _17379_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24593__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19118_ _19117_/Y _19114_/X _19095_/X _19114_/X VGND VGND VPWR VPWR _23448_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11710__A _13053_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20390_ _17182_/B _20390_/B _20373_/X VGND VGND VPWR VPWR _20390_/X sky130_fd_sc_hd__and3_4
XANTENNA__24522__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15312__A1_N _13613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19049_ _19034_/Y VGND VGND VPWR VPWR _19049_/X sky130_fd_sc_hd__buf_2
XFILLER_12_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12706__B1 _12674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22060_ _21667_/X _19486_/Y VGND VGND VPWR VPWR _22060_/X sky130_fd_sc_hd__or2_4
XFILLER_82_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21011_ _21007_/X _21010_/X _24745_/Q VGND VGND VPWR VPWR _21011_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_59_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21854__A _21051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15671__A2 _15647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21573__B _21860_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22962_ _22539_/X _22960_/X _20750_/X _22961_/X VGND VGND VPWR VPWR _22963_/A sky130_fd_sc_hd__o22a_4
XANTENNA__22941__B2 _22029_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24701_ _24698_/CLK _24701_/D HRESETn VGND VGND VPWR VPWR _24701_/Q sky130_fd_sc_hd__dfrtp_4
X_21913_ _21913_/A _21913_/B VGND VGND VPWR VPWR _21914_/C sky130_fd_sc_hd__or2_4
XFILLER_71_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22893_ _22163_/A _22892_/X VGND VGND VPWR VPWR _22893_/X sky130_fd_sc_hd__and2_4
XANTENNA__15423__A2 _15415_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24632_ _23618_/CLK _15273_/X HRESETn VGND VGND VPWR VPWR _15270_/A sky130_fd_sc_hd__dfstp_4
X_21844_ _21843_/X VGND VGND VPWR VPWR _21844_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21775_ _21764_/A _21773_/X _21774_/X VGND VGND VPWR VPWR _21775_/X sky130_fd_sc_hd__and3_4
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24563_ _25123_/CLK _24563_/D HRESETn VGND VGND VPWR VPWR _12117_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20726_ _24026_/Q _24024_/Q _24025_/Q _20725_/X VGND VGND VPWR VPWR _20726_/X sky130_fd_sc_hd__o22a_4
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23514_ _23514_/CLK _23514_/D VGND VGND VPWR VPWR _17870_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_51_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16384__B1 _16291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24494_ _25090_/CLK _24494_/D HRESETn VGND VGND VPWR VPWR _24494_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_213_0_HCLK clkbuf_8_213_0_HCLK/A VGND VGND VPWR VPWR _23824_/CLK sky130_fd_sc_hd__clkbuf_1
X_20657_ _20656_/Y _20653_/Y _20660_/B VGND VGND VPWR VPWR _20657_/X sky130_fd_sc_hd__o21a_4
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23445_ _23469_/CLK _23445_/D VGND VGND VPWR VPWR _17714_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19322__B1 _19207_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11620__A _13668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23376_ _23471_/CLK _23376_/D VGND VGND VPWR VPWR _13277_/B sky130_fd_sc_hd__dfxtp_4
X_20588_ _16537_/Y _20574_/X _20583_/X _20587_/X VGND VGND VPWR VPWR _20589_/A sky130_fd_sc_hd__o22a_4
XANTENNA__24263__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22209__B1 _11532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12861__A2_N _24459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25115_ _25115_/CLK _12261_/X HRESETn VGND VGND VPWR VPWR _25115_/Q sky130_fd_sc_hd__dfrtp_4
X_22327_ _20605_/Y _22279_/X _20468_/Y _20926_/X VGND VGND VPWR VPWR _22327_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16687__B2 _17482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23666__D _23666_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13060_ _23890_/Q VGND VGND VPWR VPWR _13297_/A sky130_fd_sc_hd__buf_2
X_22258_ _22258_/A _22299_/A VGND VGND VPWR VPWR _22258_/X sky130_fd_sc_hd__and2_4
X_25046_ _25046_/CLK _12749_/X HRESETn VGND VGND VPWR VPWR _12581_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24870__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12011_ _12011_/A VGND VGND VPWR VPWR _12011_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21209_ _21374_/A _21209_/B VGND VGND VPWR VPWR _21209_/X sky130_fd_sc_hd__or2_4
XANTENNA__21725__A1_N _11999_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22189_ _22444_/B _22187_/X _21046_/X _12582_/A _22188_/X VGND VGND VPWR VPWR _22189_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12451__A _12451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16858__A _16858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15662__A2 _15647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16750_ _20737_/B _16748_/X _16749_/Y VGND VGND VPWR VPWR _16750_/X sky130_fd_sc_hd__o21a_4
XFILLER_115_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13962_ _24892_/Q _13930_/B _24892_/Q _13930_/B VGND VGND VPWR VPWR _13962_/X sky130_fd_sc_hd__a2bb2o_4
X_15701_ _12307_/Y _15698_/X _15390_/X _15698_/X VGND VGND VPWR VPWR _15701_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12913_ _12922_/A _12908_/B _12913_/C VGND VGND VPWR VPWR _12914_/A sky130_fd_sc_hd__or3_4
XANTENNA__22932__B2 _22531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25051__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16681_ _20919_/A _13480_/B _13463_/A _16680_/X VGND VGND VPWR VPWR _16681_/X sky130_fd_sc_hd__o22a_4
X_13893_ _13886_/X VGND VGND VPWR VPWR _13893_/X sky130_fd_sc_hd__buf_2
XFILLER_94_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18420_ _18420_/A VGND VGND VPWR VPWR _18420_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13282__A _13065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15632_ _15619_/X _15617_/X _15522_/X _24505_/Q _15585_/A VGND VGND VPWR VPWR _24505_/D
+ sky130_fd_sc_hd__a32o_4
X_12844_ _12837_/X _12844_/B _12844_/C _12844_/D VGND VGND VPWR VPWR _12844_/X sky130_fd_sc_hd__or4_4
XFILLER_74_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18351_ _23834_/Q VGND VGND VPWR VPWR _18352_/A sky130_fd_sc_hd__inv_2
X_15563_ _15556_/X VGND VGND VPWR VPWR _15563_/X sky130_fd_sc_hd__buf_2
XFILLER_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12775_ _12774_/Y _24440_/Q _12774_/Y _24440_/Q VGND VGND VPWR VPWR _12775_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_23_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _24008_/Q VGND VGND VPWR VPWR _17330_/A sky130_fd_sc_hd__inv_2
XFILLER_14_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14514_ _14510_/Y _14513_/Y _14509_/X _14513_/A VGND VGND VPWR VPWR _24750_/D sky130_fd_sc_hd__o22a_4
XPHY_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11725_/X VGND VGND VPWR VPWR _11726_/Y sky130_fd_sc_hd__inv_2
X_18282_ _18284_/A _18282_/B _18281_/Y VGND VGND VPWR VPWR _23862_/D sky130_fd_sc_hd__and3_4
XPHY_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ HWDATA[16] VGND VGND VPWR VPWR _15494_/X sky130_fd_sc_hd__buf_2
XPHY_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17233_ _11745_/B _11759_/X _17233_/C _17233_/D VGND VGND VPWR VPWR _17233_/X sky130_fd_sc_hd__or4_4
X_14445_ _14445_/A VGND VGND VPWR VPWR _14445_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22448__B1 _20780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _11657_/A VGND VGND VPWR VPWR _13559_/A sky130_fd_sc_hd__inv_2
XPHY_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11530__A _22992_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19313__B1 _19311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17164_ _17161_/A _17161_/B VGND VGND VPWR VPWR _17164_/Y sky130_fd_sc_hd__nand2_4
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14376_ _14420_/A _14420_/B VGND VGND VPWR VPWR _14377_/B sky130_fd_sc_hd__and2_4
X_11588_ _11599_/A VGND VGND VPWR VPWR _11588_/X sky130_fd_sc_hd__buf_2
XANTENNA__20843__A _11725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16115_ _21716_/A _16112_/X _15897_/X _16112_/X VGND VGND VPWR VPWR _24329_/D sky130_fd_sc_hd__a2bb2o_4
X_13327_ _16301_/A _21707_/B VGND VGND VPWR VPWR _13328_/A sky130_fd_sc_hd__or2_4
X_17095_ _17040_/A _17116_/A _17116_/B VGND VGND VPWR VPWR _17096_/B sky130_fd_sc_hd__or3_4
XANTENNA__19409__A _19396_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16046_ _16046_/A VGND VGND VPWR VPWR _16046_/X sky130_fd_sc_hd__buf_2
X_13258_ _11732_/B _13258_/B VGND VGND VPWR VPWR _13258_/X sky130_fd_sc_hd__or2_4
XFILLER_83_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23986__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12209_ _12209_/A VGND VGND VPWR VPWR _12214_/B sky130_fd_sc_hd__inv_2
XANTENNA__21423__B2 _22610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13189_ _13221_/A _13189_/B _13189_/C VGND VGND VPWR VPWR _13190_/C sky130_fd_sc_hd__and3_4
XFILLER_123_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23915__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19805_ _19800_/X _18067_/X _13668_/A _23204_/Q _19802_/X VGND VGND VPWR VPWR _19805_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_111_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25139__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17997_ _11671_/Y _17995_/X _17205_/X _17995_/X VGND VGND VPWR VPWR _17997_/X sky130_fd_sc_hd__a2bb2o_4
X_16948_ _16778_/Y _16952_/B VGND VGND VPWR VPWR _16953_/A sky130_fd_sc_hd__or2_4
X_19736_ _19531_/A _18038_/X _23903_/Q _18031_/B VGND VGND VPWR VPWR _19737_/A sky130_fd_sc_hd__or4_4
XFILLER_133_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_105_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_211_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16879_ _16879_/A _17067_/A VGND VGND VPWR VPWR _16879_/X sky130_fd_sc_hd__and2_4
X_19667_ _19667_/A VGND VGND VPWR VPWR _19680_/A sky130_fd_sc_hd__inv_2
XFILLER_42_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18618_ _23640_/Q _18617_/X VGND VGND VPWR VPWR _18619_/B sky130_fd_sc_hd__or2_4
X_19598_ _19594_/Y _19596_/X _19597_/X _19596_/X VGND VGND VPWR VPWR _23278_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17599__A _16700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18549_ _18548_/X VGND VGND VPWR VPWR _23817_/D sky130_fd_sc_hd__inv_2
XANTENNA__24774__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21560_ _22943_/A _21548_/X _21559_/Y VGND VGND VPWR VPWR _21706_/A sky130_fd_sc_hd__o21ai_4
XFILLER_33_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24703__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20511_ _20511_/A VGND VGND VPWR VPWR _20511_/X sky130_fd_sc_hd__buf_2
XFILLER_21_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21491_ _21491_/A _21490_/X VGND VGND VPWR VPWR _21496_/B sky130_fd_sc_hd__or2_4
XFILLER_14_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22952__B _22952_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23230_ _23246_/CLK _23230_/D VGND VGND VPWR VPWR _23230_/Q sky130_fd_sc_hd__dfxtp_4
X_20442_ _13506_/B VGND VGND VPWR VPWR _20442_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16118__B1 _15992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20753__A _20753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14965__A2_N _24258_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23161_ _25112_/CLK _19919_/X VGND VGND VPWR VPWR _19917_/A sky130_fd_sc_hd__dfxtp_4
X_20373_ _17187_/A VGND VGND VPWR VPWR _20373_/X sky130_fd_sc_hd__buf_2
XFILLER_101_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_43_0_HCLK clkbuf_8_43_0_HCLK/A VGND VGND VPWR VPWR _23563_/CLK sky130_fd_sc_hd__clkbuf_1
X_22112_ _20968_/X _22108_/X _22111_/X VGND VGND VPWR VPWR _22112_/X sky130_fd_sc_hd__or3_4
XANTENNA__14144__A2 _23042_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23092_ _23100_/CLK _20101_/X VGND VGND VPWR VPWR _23092_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13352__B1 _11636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12155__B2 _24575_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22043_ _22043_/A _21638_/X VGND VGND VPWR VPWR _22043_/X sky130_fd_sc_hd__or2_4
XFILLER_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23656__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16678__A _17725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23994_ _25214_/CLK _17392_/X HRESETn VGND VGND VPWR VPWR _17309_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22914__A1 _23026_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21717__A2 _21716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22914__B2 _22460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22945_ _16400_/Y _21715_/X _14740_/Y _22225_/A VGND VGND VPWR VPWR _22945_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17200__A2_N _17198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11615__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22876_ _14714_/A _22745_/B VGND VGND VPWR VPWR _22876_/X sky130_fd_sc_hd__or2_4
XFILLER_44_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20928__A _20900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24615_ _23734_/CLK _15323_/X HRESETn VGND VGND VPWR VPWR _23026_/A sky130_fd_sc_hd__dfrtp_4
X_21827_ _21913_/A _21827_/B VGND VGND VPWR VPWR _21827_/X sky130_fd_sc_hd__or2_4
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14926__A _24257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ _24529_/Q VGND VGND VPWR VPWR _12560_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16357__B1 _16096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24546_ _24566_/CLK _15525_/X HRESETn VGND VGND VPWR VPWR _24546_/Q sky130_fd_sc_hd__dfrtp_4
X_21758_ _15572_/A _23034_/B VGND VGND VPWR VPWR _21758_/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24444__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11511_ _24619_/Q VGND VGND VPWR VPWR _16038_/B sky130_fd_sc_hd__inv_2
XFILLER_54_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20709_ _20709_/A VGND VGND VPWR VPWR _20710_/A sky130_fd_sc_hd__inv_2
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12491_ _12465_/B _12464_/X _12453_/X _12487_/Y VGND VGND VPWR VPWR _12492_/A sky130_fd_sc_hd__a211o_4
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24477_ _24307_/CLK _15696_/X HRESETn VGND VGND VPWR VPWR _24477_/Q sky130_fd_sc_hd__dfrtp_4
X_21689_ _20782_/X _21672_/X _21688_/X VGND VGND VPWR VPWR _21689_/X sky130_fd_sc_hd__and3_4
XFILLER_71_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14230_ _14230_/A VGND VGND VPWR VPWR _14230_/Y sky130_fd_sc_hd__inv_2
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23428_ _25067_/CLK _19176_/X VGND VGND VPWR VPWR _19174_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14161_ _14160_/X VGND VGND VPWR VPWR _14161_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21478__B _19656_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23359_ _24998_/CLK _23359_/D VGND VGND VPWR VPWR _13306_/B sky130_fd_sc_hd__dfxtp_4
X_13112_ _13026_/X _13107_/X _13112_/C VGND VGND VPWR VPWR _13113_/C sky130_fd_sc_hd__or3_4
XANTENNA__14135__A2 _14122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14092_ _14090_/Y _14091_/X _13638_/X _14091_/X VGND VGND VPWR VPWR _24857_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13277__A _13309_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13043_ _13047_/A _13043_/B _13043_/C VGND VGND VPWR VPWR _13043_/X sky130_fd_sc_hd__and3_4
X_17920_ _17821_/A _17920_/B VGND VGND VPWR VPWR _17920_/X sky130_fd_sc_hd__or2_4
X_25029_ _24432_/CLK _12924_/Y HRESETn VGND VGND VPWR VPWR _22778_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17851_ _17947_/A _17851_/B _17851_/C VGND VGND VPWR VPWR _17851_/X sky130_fd_sc_hd__or3_4
XFILLER_65_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16802_ _24081_/Q VGND VGND VPWR VPWR _16802_/Y sky130_fd_sc_hd__inv_2
X_17782_ _17782_/A _17782_/B VGND VGND VPWR VPWR _17783_/C sky130_fd_sc_hd__or2_4
X_14994_ _14994_/A VGND VGND VPWR VPWR _24710_/D sky130_fd_sc_hd__inv_2
XANTENNA__21708__A2 _11954_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22905__A1 _22201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16733_ _22920_/A VGND VGND VPWR VPWR _16733_/Y sky130_fd_sc_hd__inv_2
X_19521_ _21517_/B _19516_/X _19455_/X _19516_/X VGND VGND VPWR VPWR _23306_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13945_ _13944_/X VGND VGND VPWR VPWR _13945_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20916__B1 _13441_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19452_ _19452_/A VGND VGND VPWR VPWR _19452_/X sky130_fd_sc_hd__buf_2
XANTENNA__11525__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16664_ _14726_/Y _16663_/X _16455_/X _16663_/X VGND VGND VPWR VPWR _16664_/X sky130_fd_sc_hd__a2bb2o_4
X_13876_ _13833_/A _13880_/B _13828_/D _13876_/D VGND VGND VPWR VPWR _13877_/D sky130_fd_sc_hd__and4_4
XANTENNA__16596__B1 _15497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15615_ _15611_/X _15599_/X _15499_/X _24516_/Q _15612_/X VGND VGND VPWR VPWR _24516_/D
+ sky130_fd_sc_hd__a32o_4
X_18403_ _16398_/Y _23843_/Q _16398_/Y _23843_/Q VGND VGND VPWR VPWR _18403_/X sky130_fd_sc_hd__a2bb2o_4
X_12827_ _21851_/A VGND VGND VPWR VPWR _12827_/Y sky130_fd_sc_hd__inv_2
X_19383_ _13216_/B VGND VGND VPWR VPWR _19383_/Y sky130_fd_sc_hd__inv_2
X_16595_ _16584_/A VGND VGND VPWR VPWR _16595_/X sky130_fd_sc_hd__buf_2
XFILLER_43_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18334_ _18334_/A _18333_/Y VGND VGND VPWR VPWR _18335_/B sky130_fd_sc_hd__or2_4
XFILLER_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15546_ _15558_/A VGND VGND VPWR VPWR _15546_/X sky130_fd_sc_hd__buf_2
XFILLER_37_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12758_ _12593_/A _12758_/B VGND VGND VPWR VPWR _12759_/B sky130_fd_sc_hd__or2_4
XFILLER_37_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16348__B1 _16179_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24185__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ _11708_/X VGND VGND VPWR VPWR _13053_/C sky130_fd_sc_hd__inv_2
X_18265_ _18207_/B _18265_/B VGND VGND VPWR VPWR _18268_/B sky130_fd_sc_hd__or2_4
X_15477_ HWDATA[26] VGND VGND VPWR VPWR _15477_/X sky130_fd_sc_hd__buf_2
XANTENNA__21892__B2 _21868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24114__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12689_ _12550_/X _12691_/B _12688_/Y VGND VGND VPWR VPWR _12689_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12356__A _12356_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17216_ _17215_/Y _17213_/X _16617_/X _17213_/X VGND VGND VPWR VPWR _24013_/D sky130_fd_sc_hd__a2bb2o_4
X_14428_ _14428_/A VGND VGND VPWR VPWR _21534_/A sky130_fd_sc_hd__inv_2
XFILLER_128_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18196_ _18262_/A VGND VGND VPWR VPWR _18226_/A sky130_fd_sc_hd__buf_2
XANTENNA__17985__A1_N _11691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20873__A1_N _14264_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17147_ _17034_/A _17145_/X _17146_/Y VGND VGND VPWR VPWR _24036_/D sky130_fd_sc_hd__o21a_4
X_14359_ _14352_/A _13877_/D _14359_/C _13898_/A VGND VGND VPWR VPWR _14360_/B sky130_fd_sc_hd__or4_4
XANTENNA__22841__B1 _25216_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_2_0_HCLK clkbuf_7_1_0_HCLK/X VGND VGND VPWR VPWR _23388_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__14571__A _17742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15323__A1 _11533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17078_ _17026_/B _17077_/X VGND VGND VPWR VPWR _17079_/A sky130_fd_sc_hd__or2_4
XFILLER_48_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16029_ _14564_/X _14558_/X _14560_/Y VGND VGND VPWR VPWR _16033_/B sky130_fd_sc_hd__o21a_4
XFILLER_97_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22899__A2_N _22896_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14834__B1 _14712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22012__B _20866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19719_ _21808_/B _19710_/X _19717_/X _19718_/X VGND VGND VPWR VPWR _19719_/X sky130_fd_sc_hd__a2bb2o_4
X_20991_ _14528_/A _20991_/B _20990_/X VGND VGND VPWR VPWR _20991_/X sky130_fd_sc_hd__and3_4
XANTENNA__24955__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22730_ _22730_/A _22730_/B VGND VGND VPWR VPWR _22744_/C sky130_fd_sc_hd__nor2_4
XFILLER_26_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20748__A _20747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22661_ _22661_/A _22627_/X _22661_/C _22660_/X VGND VGND VPWR VPWR HRDATA[19] sky130_fd_sc_hd__or4_4
XFILLER_55_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24400_ _24399_/CLK _15898_/X HRESETn VGND VGND VPWR VPWR _24400_/Q sky130_fd_sc_hd__dfrtp_4
X_21612_ _21612_/A _20084_/Y VGND VGND VPWR VPWR _21614_/B sky130_fd_sc_hd__or2_4
XFILLER_107_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22592_ _22116_/X _22591_/X _21974_/X _12117_/A _22118_/X VGND VGND VPWR VPWR _22592_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_107_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14274__A2_N _14268_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17000__B2 _24040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24331_ _23852_/CLK _16110_/X HRESETn VGND VGND VPWR VPWR _24331_/Q sky130_fd_sc_hd__dfrtp_4
X_21543_ _21543_/A VGND VGND VPWR VPWR _21544_/A sky130_fd_sc_hd__buf_2
XANTENNA__21883__B2 _21570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21474_ _21340_/A _21474_/B VGND VGND VPWR VPWR _21474_/X sky130_fd_sc_hd__or2_4
X_24262_ _24262_/CLK _16284_/X HRESETn VGND VGND VPWR VPWR _24262_/Q sky130_fd_sc_hd__dfrtp_4
X_20425_ _20425_/A VGND VGND VPWR VPWR _20425_/X sky130_fd_sc_hd__buf_2
XFILLER_101_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23213_ _23282_/CLK _19784_/X VGND VGND VPWR VPWR _19783_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_119_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24193_ _24192_/CLK _16468_/X HRESETn VGND VGND VPWR VPWR _16467_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_135_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23837__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20356_ _20355_/X VGND VGND VPWR VPWR _23669_/D sky130_fd_sc_hd__inv_2
X_23144_ _25044_/CLK _23144_/D VGND VGND VPWR VPWR _23144_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12128__B2 _24557_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23075_ _23993_/CLK _20139_/X VGND VGND VPWR VPWR _23075_/Q sky130_fd_sc_hd__dfxtp_4
X_20287_ _20286_/X VGND VGND VPWR VPWR _20287_/X sky130_fd_sc_hd__buf_2
XFILLER_122_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16502__A1_N _16501_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22026_ _14286_/Y _12063_/X _20331_/A _22227_/B VGND VGND VPWR VPWR _22026_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20071__B1 _19963_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14842__A2_N _24148_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11639__B1 _25191_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22899__B1 _22677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11991_ _11985_/Y _11990_/X _11604_/X _11990_/X VGND VGND VPWR VPWR _25147_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24696__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23977_ _24962_/CLK _17469_/X HRESETn VGND VGND VPWR VPWR _17466_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_17_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22857__B _22857_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13730_ _13730_/A VGND VGND VPWR VPWR _13730_/X sky130_fd_sc_hd__buf_2
XFILLER_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22928_ _24218_/Q _23020_/B VGND VGND VPWR VPWR _22928_/X sky130_fd_sc_hd__or2_4
XANTENNA__16578__B1 _16153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14857__A2_N _24156_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13661_ _13647_/Y VGND VGND VPWR VPWR _13661_/X sky130_fd_sc_hd__buf_2
XFILLER_73_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22859_ _22859_/A VGND VGND VPWR VPWR _22859_/X sky130_fd_sc_hd__buf_2
XANTENNA__20042__A2_N _20036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15400_ _24586_/Q VGND VGND VPWR VPWR _21285_/A sky130_fd_sc_hd__inv_2
X_12612_ _25059_/Q VGND VGND VPWR VPWR _12612_/Y sky130_fd_sc_hd__inv_2
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16380_ _16378_/Y _16372_/X _15992_/X _16379_/X VGND VGND VPWR VPWR _24226_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13592_ _13561_/B _13580_/X _13591_/Y _13587_/X _24954_/Q VGND VGND VPWR VPWR _24954_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15331_ _15331_/A VGND VGND VPWR VPWR _15331_/Y sky130_fd_sc_hd__inv_2
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12543_ _12649_/C _24513_/Q _12649_/C _24513_/Q VGND VGND VPWR VPWR _12543_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24529_ _25005_/CLK _15594_/X HRESETn VGND VGND VPWR VPWR _24529_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18050_ _18049_/X _18036_/X _18049_/X _18036_/X VGND VGND VPWR VPWR _18050_/X sky130_fd_sc_hd__a2bb2o_4
X_15262_ _15262_/A VGND VGND VPWR VPWR _15262_/X sky130_fd_sc_hd__buf_2
XANTENNA__22977__A1_N _21546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12474_ _12412_/A _12412_/B _12474_/C _12466_/B VGND VGND VPWR VPWR _12480_/B sky130_fd_sc_hd__or4_4
X_17001_ _16160_/Y _17089_/A _16160_/Y _17089_/A VGND VGND VPWR VPWR _17001_/X sky130_fd_sc_hd__a2bb2o_4
X_14213_ _15801_/A VGND VGND VPWR VPWR _14213_/X sky130_fd_sc_hd__buf_2
XFILLER_125_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15193_ _14939_/Y _15188_/B _15190_/B _15147_/X VGND VGND VPWR VPWR _15193_/X sky130_fd_sc_hd__a211o_4
XFILLER_126_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14144_ _20889_/A _23042_/B _24839_/Q VGND VGND VPWR VPWR _24840_/D sky130_fd_sc_hd__a21o_4
XFILLER_10_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16502__B1 _16254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14075_ _23689_/Q _14071_/X _14074_/X VGND VGND VPWR VPWR _14075_/Y sky130_fd_sc_hd__a21oi_4
X_18952_ _17839_/B VGND VGND VPWR VPWR _18952_/Y sky130_fd_sc_hd__inv_2
X_13026_ _13271_/A VGND VGND VPWR VPWR _13026_/X sky130_fd_sc_hd__buf_2
X_17903_ _17903_/A _17903_/B VGND VGND VPWR VPWR _17903_/X sky130_fd_sc_hd__or2_4
X_18883_ _18743_/X VGND VGND VPWR VPWR _18883_/X sky130_fd_sc_hd__buf_2
XANTENNA__22113__A _21339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17834_ _17796_/X _17834_/B VGND VGND VPWR VPWR _17834_/X sky130_fd_sc_hd__or2_4
XFILLER_66_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14977_ _14987_/A _15094_/A _14977_/C _14990_/A VGND VGND VPWR VPWR _14980_/B sky130_fd_sc_hd__or4_4
X_17765_ _15728_/A VGND VGND VPWR VPWR _17765_/X sky130_fd_sc_hd__buf_2
XFILLER_81_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19504_ _21197_/B _19501_/X _19462_/X _19501_/X VGND VGND VPWR VPWR _23312_/D sky130_fd_sc_hd__a2bb2o_4
X_13928_ _24888_/Q _13928_/B _13928_/C VGND VGND VPWR VPWR _13928_/X sky130_fd_sc_hd__or3_4
X_16716_ _16709_/X _16716_/B _16716_/C _16716_/D VGND VGND VPWR VPWR _16716_/X sky130_fd_sc_hd__or4_4
X_17696_ _17692_/X _17695_/X _16678_/X VGND VGND VPWR VPWR _17696_/X sky130_fd_sc_hd__o21a_4
XFILLER_35_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24366__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16647_ _16627_/A VGND VGND VPWR VPWR _16647_/X sky130_fd_sc_hd__buf_2
X_19435_ _19434_/Y _19432_/X _19366_/X _19432_/X VGND VGND VPWR VPWR _23336_/D sky130_fd_sc_hd__a2bb2o_4
X_13859_ _13815_/X VGND VGND VPWR VPWR _13861_/A sky130_fd_sc_hd__inv_2
XANTENNA__19290__A2_N _19284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16578_ _14859_/Y _16576_/X _16153_/X _16576_/X VGND VGND VPWR VPWR _24151_/D sky130_fd_sc_hd__a2bb2o_4
X_19366_ _18801_/X VGND VGND VPWR VPWR _19366_/X sky130_fd_sc_hd__buf_2
XANTENNA__22783__A _22783_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15529_ _15422_/A _15531_/B VGND VGND VPWR VPWR _15529_/X sky130_fd_sc_hd__or2_4
X_18317_ _18290_/X _18304_/X _18317_/C VGND VGND VPWR VPWR _18317_/X sky130_fd_sc_hd__and3_4
X_19297_ _21352_/B _19296_/X _11857_/X _19296_/X VGND VGND VPWR VPWR _19297_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18248_ _18559_/B _18248_/B _18248_/C VGND VGND VPWR VPWR _18249_/A sky130_fd_sc_hd__or3_4
XFILLER_129_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18179_ _23873_/Q VGND VGND VPWR VPWR _18179_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20210_ _20209_/X VGND VGND VPWR VPWR _20210_/X sky130_fd_sc_hd__buf_2
XANTENNA__23930__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21190_ _21189_/X VGND VGND VPWR VPWR _21190_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25154__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20141_ _20141_/A VGND VGND VPWR VPWR _20141_/X sky130_fd_sc_hd__buf_2
XFILLER_131_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14935__A1_N _24667_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_117_0_HCLK clkbuf_7_58_0_HCLK/X VGND VGND VPWR VPWR _23661_/CLK sky130_fd_sc_hd__clkbuf_1
X_20072_ _20072_/A VGND VGND VPWR VPWR _20072_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13645__A _14218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19994__B1 _19421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23900_ _23343_/CLK _18041_/X HRESETn VGND VGND VPWR VPWR _18022_/A sky130_fd_sc_hd__dfrtp_4
X_24880_ _23648_/CLK _24880_/D HRESETn VGND VGND VPWR VPWR _13925_/C sky130_fd_sc_hd__dfrtp_4
X_23831_ _24654_/CLK _23831_/D HRESETn VGND VGND VPWR VPWR _23831_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23625__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15480__B1 _24570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23762_ _23762_/CLK _23762_/D HRESETn VGND VGND VPWR VPWR HREADYOUT sky130_fd_sc_hd__dfstp_4
X_20974_ _20979_/A _20974_/B VGND VGND VPWR VPWR _20974_/X sky130_fd_sc_hd__or2_4
XFILLER_53_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20765__A1_N _21357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22713_ _12410_/Y _22606_/X _24048_/Q _22652_/X VGND VGND VPWR VPWR _22716_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14476__A _14429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24036__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23693_ _24897_/CLK _20237_/X HRESETn VGND VGND VPWR VPWR _23693_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15232__B1 _15126_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22644_ _22249_/A VGND VGND VPWR VPWR _22897_/B sky130_fd_sc_hd__buf_2
XFILLER_15_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22575_ _22840_/A VGND VGND VPWR VPWR _22576_/A sky130_fd_sc_hd__buf_2
XFILLER_51_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24314_ _24037_/CLK _16156_/X HRESETn VGND VGND VPWR VPWR _24314_/Q sky130_fd_sc_hd__dfrtp_4
X_21526_ _21500_/A _21524_/X _21525_/X VGND VGND VPWR VPWR _21526_/X sky130_fd_sc_hd__and3_4
X_24245_ _24213_/CLK _16329_/X HRESETn VGND VGND VPWR VPWR _24245_/Q sky130_fd_sc_hd__dfrtp_4
X_21457_ _21457_/A _21457_/B _21457_/C _21457_/D VGND VGND VPWR VPWR _21457_/X sky130_fd_sc_hd__or4_4
XANTENNA__13010__A2 _12921_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23671__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15100__A _15159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12190_ _12190_/A _12190_/B _12190_/C VGND VGND VPWR VPWR _12190_/X sky130_fd_sc_hd__and3_4
X_20408_ _20203_/Y _20264_/A _20202_/Y VGND VGND VPWR VPWR _20409_/C sky130_fd_sc_hd__o21a_4
X_21388_ _21384_/X _21387_/X _21231_/X VGND VGND VPWR VPWR _21396_/B sky130_fd_sc_hd__o21a_4
XFILLER_135_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24176_ _24177_/CLK _16512_/X HRESETn VGND VGND VPWR VPWR _24176_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_13_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_134_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23127_ _23128_/CLK _23127_/D VGND VGND VPWR VPWR _20007_/A sky130_fd_sc_hd__dfxtp_4
X_20339_ _20183_/X _20191_/B _13916_/X VGND VGND VPWR VPWR _23650_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_7_76_0_HCLK clkbuf_7_76_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_76_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23058_ _20736_/X VGND VGND VPWR VPWR IRQ[6] sky130_fd_sc_hd__buf_2
XANTENNA__24877__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14900_ _14900_/A VGND VGND VPWR VPWR _14900_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19985__B1 _15561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22009_ _20447_/Y _20819_/X _22584_/A _22008_/X VGND VGND VPWR VPWR _22009_/X sky130_fd_sc_hd__o22a_4
XFILLER_27_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17027__A _17027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15880_ _15885_/A VGND VGND VPWR VPWR _15880_/X sky130_fd_sc_hd__buf_2
XANTENNA__16799__B1 _24423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21792__B1 _21642_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14831_ _14831_/A VGND VGND VPWR VPWR _14831_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22587__B _22587_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17550_ _17499_/X _17550_/B VGND VGND VPWR VPWR _17550_/X sky130_fd_sc_hd__or2_4
XANTENNA__15770__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14762_ _24695_/Q VGND VGND VPWR VPWR _14762_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21491__B _21490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11974_ _11973_/Y _11971_/X _11626_/X _11971_/X VGND VGND VPWR VPWR _25152_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18004__A3 _16558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16501_ _24180_/Q VGND VGND VPWR VPWR _16501_/Y sky130_fd_sc_hd__inv_2
X_13713_ _23685_/Q VGND VGND VPWR VPWR _13794_/A sky130_fd_sc_hd__buf_2
XFILLER_45_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17481_ _17481_/A VGND VGND VPWR VPWR _17481_/Y sky130_fd_sc_hd__inv_2
X_14693_ pwm_S6 VGND VGND VPWR VPWR _14693_/Y sky130_fd_sc_hd__inv_2
X_16432_ _24206_/Q VGND VGND VPWR VPWR _16432_/Y sky130_fd_sc_hd__inv_2
X_19220_ _23411_/Q VGND VGND VPWR VPWR _19220_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13644_ _13644_/A VGND VGND VPWR VPWR _14218_/A sky130_fd_sc_hd__buf_2
XFILLER_71_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19151_ _23436_/Q VGND VGND VPWR VPWR _19151_/Y sky130_fd_sc_hd__inv_2
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16363_ _16363_/A VGND VGND VPWR VPWR _16363_/Y sky130_fd_sc_hd__inv_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _13572_/A _13571_/X VGND VGND VPWR VPWR _13575_/Y sky130_fd_sc_hd__nand2_4
XFILLER_73_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18102_ _18101_/X VGND VGND VPWR VPWR _18102_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23759__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15314_ _15314_/A _15314_/B VGND VGND VPWR VPWR _15314_/X sky130_fd_sc_hd__or2_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12526_ _12456_/X _12505_/B _12526_/C VGND VGND VPWR VPWR _12526_/X sky130_fd_sc_hd__and3_4
X_19082_ _19081_/Y _19079_/X _19038_/X _19079_/X VGND VGND VPWR VPWR _23461_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16294_ _24255_/Q VGND VGND VPWR VPWR _16294_/Y sky130_fd_sc_hd__inv_2
X_18033_ _23901_/Q _18022_/A VGND VGND VPWR VPWR _18033_/X sky130_fd_sc_hd__and2_4
X_15245_ _15251_/B VGND VGND VPWR VPWR _15245_/X sky130_fd_sc_hd__buf_2
X_12457_ _12456_/X VGND VGND VPWR VPWR _12460_/A sky130_fd_sc_hd__buf_2
XANTENNA__12634__A _12933_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15176_ _15165_/A _15170_/X _15176_/C VGND VGND VPWR VPWR _24668_/D sky130_fd_sc_hd__and3_4
XANTENNA__21947__A _21393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12388_ _25073_/Q VGND VGND VPWR VPWR _12388_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14127_ _14115_/X VGND VGND VPWR VPWR _14127_/X sky130_fd_sc_hd__buf_2
X_19984_ _23136_/Q VGND VGND VPWR VPWR _21233_/B sky130_fd_sc_hd__inv_2
XFILLER_125_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14058_ _14057_/Y _14053_/X _13635_/X _14053_/X VGND VGND VPWR VPWR _14058_/X sky130_fd_sc_hd__a2bb2o_4
X_18935_ _18935_/A VGND VGND VPWR VPWR _18935_/X sky130_fd_sc_hd__buf_2
XFILLER_97_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14501__A2 _14480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12512__A1 _12406_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13009_ _13009_/A VGND VGND VPWR VPWR _13009_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19976__B1 _19448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18866_ _18854_/A VGND VGND VPWR VPWR _18866_/X sky130_fd_sc_hd__buf_2
XFILLER_121_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24547__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17817_ _17817_/A _19177_/A VGND VGND VPWR VPWR _17818_/C sky130_fd_sc_hd__or2_4
XFILLER_39_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18797_ _23561_/Q VGND VGND VPWR VPWR _18797_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22327__A2 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22497__B _22497_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19152__A _18743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17748_ _17895_/A _19081_/A VGND VGND VPWR VPWR _17751_/B sky130_fd_sc_hd__or2_4
XANTENNA__21535__B1 _21256_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17203__B2 _17198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17679_ _17676_/X _17679_/B _17679_/C VGND VGND VPWR VPWR _17679_/X sky130_fd_sc_hd__and3_4
XFILLER_1_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19418_ _19417_/Y VGND VGND VPWR VPWR _19418_/X sky130_fd_sc_hd__buf_2
X_20690_ _11886_/X _20691_/B VGND VGND VPWR VPWR _20690_/X sky130_fd_sc_hd__and2_4
XFILLER_91_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19349_ _19349_/A VGND VGND VPWR VPWR _19349_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19900__B1 _19835_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22360_ _21642_/X VGND VGND VPWR VPWR _22360_/X sky130_fd_sc_hd__buf_2
XANTENNA__22018__A _14916_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21311_ _14259_/Y _11503_/A _24786_/Q _20759_/X VGND VGND VPWR VPWR _21311_/X sky130_fd_sc_hd__a2bb2o_4
X_22291_ _22291_/A VGND VGND VPWR VPWR _22292_/D sky130_fd_sc_hd__inv_2
X_21242_ _14440_/X VGND VGND VPWR VPWR _21242_/X sky130_fd_sc_hd__buf_2
X_24030_ _24289_/CLK _17163_/X HRESETn VGND VGND VPWR VPWR _24030_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20761__A _21448_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21173_ _21167_/X _21171_/X _21172_/X VGND VGND VPWR VPWR _21174_/C sky130_fd_sc_hd__o21a_4
XANTENNA__15855__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20124_ _20122_/Y _20123_/Y _15520_/X _20123_/Y VGND VGND VPWR VPWR _23082_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24970__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20055_ _17979_/X _14197_/A VGND VGND VPWR VPWR _20055_/X sky130_fd_sc_hd__or2_4
X_24932_ _24974_/CLK _13664_/X HRESETn VGND VGND VPWR VPWR _24932_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24288__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22688__A _24114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12599__A2_N _24514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24863_ _24643_/CLK _14076_/X HRESETn VGND VGND VPWR VPWR sda_oen_o_S5 sky130_fd_sc_hd__dfstp_4
XFILLER_133_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24217__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23814_ _23824_/CLK _18558_/X HRESETn VGND VGND VPWR VPWR _23814_/Q sky130_fd_sc_hd__dfrtp_4
X_24794_ _24776_/CLK _14281_/X HRESETn VGND VGND VPWR VPWR _24794_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_38_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ _24177_/CLK _23745_/D HRESETn VGND VGND VPWR VPWR _20635_/B sky130_fd_sc_hd__dfrtp_4
X_20957_ _20971_/A VGND VGND VPWR VPWR _20964_/A sky130_fd_sc_hd__buf_2
XPHY_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _13566_/C VGND VGND VPWR VPWR _13572_/A sky130_fd_sc_hd__inv_2
XPHY_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23676_ _23676_/CLK _20388_/Y HRESETn VGND VGND VPWR VPWR _20385_/A sky130_fd_sc_hd__dfrtp_4
X_20888_ _20872_/X _20886_/Y _20887_/Y _12011_/Y _11527_/Y VGND VGND VPWR VPWR _20888_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22627_ _22348_/X _22620_/X _22622_/X _22585_/X _22626_/Y VGND VGND VPWR VPWR _22627_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23852__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13360_ _13360_/A VGND VGND VPWR VPWR _22745_/B sky130_fd_sc_hd__buf_2
XANTENNA__22573__D _22572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25076__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22558_ _21107_/X VGND VGND VPWR VPWR _22558_/X sky130_fd_sc_hd__buf_2
XFILLER_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12311_ _12451_/A _24492_/Q _12451_/A _24492_/Q VGND VGND VPWR VPWR _12312_/D sky130_fd_sc_hd__a2bb2o_4
X_21509_ _21211_/A _21509_/B VGND VGND VPWR VPWR _21509_/X sky130_fd_sc_hd__or2_4
XANTENNA__25005__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13291_ _13016_/A _18870_/A VGND VGND VPWR VPWR _13292_/C sky130_fd_sc_hd__or2_4
X_22489_ _22322_/X _22487_/X _22280_/X _22488_/X VGND VGND VPWR VPWR _22490_/B sky130_fd_sc_hd__o22a_4
XANTENNA__22870__B _22870_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15030_ _15035_/A _15034_/A _15033_/A _15020_/X VGND VGND VPWR VPWR _15036_/B sky130_fd_sc_hd__or4_4
XFILLER_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12242_ _12083_/X _12252_/B VGND VGND VPWR VPWR _12243_/B sky130_fd_sc_hd__or2_4
XANTENNA__21767__A _21519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24228_ _24201_/CLK _16374_/X HRESETn VGND VGND VPWR VPWR _16371_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15765__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12173_ _12094_/Y _12083_/X _12173_/C _12237_/A VGND VGND VPWR VPWR _12173_/X sky130_fd_sc_hd__or4_4
X_24159_ _24349_/CLK _16554_/X HRESETn VGND VGND VPWR VPWR _16553_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22038__A2_N _11961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16981_ _16981_/A _16981_/B _16978_/X _16980_/X VGND VGND VPWR VPWR _16981_/X sky130_fd_sc_hd__or4_4
XANTENNA__19958__B1 _15522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18720_ _18718_/Y _18719_/X _17205_/X _18719_/X VGND VGND VPWR VPWR _23588_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_100_0_HCLK clkbuf_7_50_0_HCLK/X VGND VGND VPWR VPWR _24623_/CLK sky130_fd_sc_hd__clkbuf_1
X_15932_ _15931_/Y _15929_/X _15837_/X _15929_/X VGND VGND VPWR VPWR _15932_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22598__A _22598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24640__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_163_0_HCLK clkbuf_7_81_0_HCLK/X VGND VGND VPWR VPWR _23154_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_49_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_6_0_HCLK clkbuf_7_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_15863_ _15862_/Y _15860_/X _15775_/X _15860_/X VGND VGND VPWR VPWR _24413_/D sky130_fd_sc_hd__a2bb2o_4
X_18651_ _18649_/Y _18645_/X _15550_/X _18650_/X VGND VGND VPWR VPWR _23612_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11517__B _15916_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17984__A2 _15430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14814_ _14814_/A VGND VGND VPWR VPWR _14814_/Y sky130_fd_sc_hd__inv_2
X_17602_ _16700_/X _17605_/B VGND VGND VPWR VPWR _17602_/Y sky130_fd_sc_hd__nand2_4
XFILLER_92_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15794_ _12778_/Y _15791_/X _15390_/X _15791_/X VGND VGND VPWR VPWR _15794_/X sky130_fd_sc_hd__a2bb2o_4
X_18582_ _18582_/A _18571_/X _18576_/X _18581_/X VGND VGND VPWR VPWR _18582_/X sky130_fd_sc_hd__or4_4
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14745_ _24691_/Q _14744_/A _14743_/X _14744_/Y VGND VGND VPWR VPWR _14745_/X sky130_fd_sc_hd__o22a_4
X_17533_ _17481_/Y _17532_/X VGND VGND VPWR VPWR _17534_/B sky130_fd_sc_hd__or2_4
X_11957_ _15422_/A _11956_/X VGND VGND VPWR VPWR _11957_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__11533__A _11532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17464_ _23976_/Q _17452_/A _17463_/X VGND VGND VPWR VPWR _17465_/A sky130_fd_sc_hd__a21o_4
XANTENNA__12032__A1_N _25144_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14676_ _14609_/A _14683_/A _14681_/A _14633_/X VGND VGND VPWR VPWR _14676_/X sky130_fd_sc_hd__or4_4
X_11888_ _11882_/B VGND VGND VPWR VPWR _11888_/Y sky130_fd_sc_hd__inv_2
X_16415_ _16413_/Y _16409_/X _16251_/X _16414_/X VGND VGND VPWR VPWR _16415_/X sky130_fd_sc_hd__a2bb2o_4
X_19203_ _23417_/Q VGND VGND VPWR VPWR _19203_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13627_ _21448_/B VGND VGND VPWR VPWR _22018_/B sky130_fd_sc_hd__buf_2
X_17395_ _17390_/A _17382_/D _17394_/X VGND VGND VPWR VPWR _23993_/D sky130_fd_sc_hd__and3_4
XFILLER_20_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16346_ _16313_/A VGND VGND VPWR VPWR _16364_/A sky130_fd_sc_hd__buf_2
X_19134_ _17846_/B VGND VGND VPWR VPWR _19134_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17220__A _13613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13558_ _13558_/A _13558_/B VGND VGND VPWR VPWR _13559_/B sky130_fd_sc_hd__or2_4
X_12509_ _12509_/A _12507_/X _12508_/X VGND VGND VPWR VPWR _25081_/D sky130_fd_sc_hd__and3_4
X_19065_ _19063_/Y _19058_/X _19041_/X _19064_/X VGND VGND VPWR VPWR _23468_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16277_ _15915_/X _16276_/X _16100_/A _22312_/A _16237_/A VGND VGND VPWR VPWR _24266_/D
+ sky130_fd_sc_hd__a32o_4
X_13489_ _11916_/X _13388_/B _13391_/B VGND VGND VPWR VPWR _13490_/B sky130_fd_sc_hd__o21a_4
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15228_ _15224_/B _15228_/B _15226_/C VGND VGND VPWR VPWR _24652_/D sky130_fd_sc_hd__and3_4
X_18016_ _17979_/X _13619_/X VGND VGND VPWR VPWR _18016_/X sky130_fd_sc_hd__or2_4
XFILLER_103_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24799__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15159_ _15159_/A _15159_/B VGND VGND VPWR VPWR _15159_/X sky130_fd_sc_hd__or2_4
XANTENNA__24728__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19967_ _23142_/Q VGND VGND VPWR VPWR _19967_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20008__B1 _15416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15683__B1 _11573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22004__C _22004_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19949__B1 _17993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18918_ _18917_/Y _18913_/X _18828_/X _18899_/Y VGND VGND VPWR VPWR _18918_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11708__A _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19898_ _21382_/B _19897_/X _19832_/X _19897_/X VGND VGND VPWR VPWR _19898_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24381__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18849_ _23543_/Q VGND VGND VPWR VPWR _18849_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24310__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13923__A scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21860_ _14887_/Y _21860_/B VGND VGND VPWR VPWR _21860_/X sky130_fd_sc_hd__and2_4
X_20811_ _24545_/Q _20799_/X _20801_/X _20810_/Y VGND VGND VPWR VPWR _20811_/X sky130_fd_sc_hd__a211o_4
XFILLER_82_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21791_ _14494_/X _21768_/Y _21776_/Y _21783_/Y _21790_/Y VGND VGND VPWR VPWR _21791_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22720__A2 _20910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19610__A _19610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23530_ _23563_/CLK _23530_/D VGND VGND VPWR VPWR _23530_/Q sky130_fd_sc_hd__dfxtp_4
X_20742_ _11725_/X VGND VGND VPWR VPWR _21113_/C sky130_fd_sc_hd__buf_2
XFILLER_1_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23461_ _24733_/CLK _23461_/D VGND VGND VPWR VPWR _19081_/A sky130_fd_sc_hd__dfxtp_4
X_20673_ _23755_/Q _13541_/X _20672_/Y VGND VGND VPWR VPWR _20673_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25200_ _24405_/CLK _25200_/D HRESETn VGND VGND VPWR VPWR _25200_/Q sky130_fd_sc_hd__dfrtp_4
X_22412_ _13535_/C _22173_/X _13508_/C _22285_/X VGND VGND VPWR VPWR _22412_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__18688__B1 _16556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23392_ _23411_/CLK _19278_/X VGND VGND VPWR VPWR _23392_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_136_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25131_ _25084_/CLK _25131_/D HRESETn VGND VGND VPWR VPWR _25131_/Q sky130_fd_sc_hd__dfrtp_4
X_22343_ _22343_/A _22281_/X VGND VGND VPWR VPWR _22343_/X sky130_fd_sc_hd__and2_4
XFILLER_30_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21587__A _21300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25062_ _25050_/CLK _12689_/X HRESETn VGND VGND VPWR VPWR _25062_/Q sky130_fd_sc_hd__dfrtp_4
X_22274_ _22354_/A _22274_/B VGND VGND VPWR VPWR _22274_/Y sky130_fd_sc_hd__nor2_4
XFILLER_128_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24013_ _24013_/CLK _24013_/D HRESETn VGND VGND VPWR VPWR _17215_/A sky130_fd_sc_hd__dfrtp_4
X_21225_ _14529_/X VGND VGND VPWR VPWR _21387_/A sky130_fd_sc_hd__buf_2
XANTENNA__15585__A _15585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24469__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21156_ _17644_/A VGND VGND VPWR VPWR _21346_/A sky130_fd_sc_hd__buf_2
XANTENNA__15674__B1 _11552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20107_ _23089_/Q VGND VGND VPWR VPWR _21474_/B sky130_fd_sc_hd__inv_2
XANTENNA__11618__A _25195_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21087_ _14093_/Y _20885_/X _24915_/Q _21720_/B VGND VGND VPWR VPWR _21087_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21747__B1 _21582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20038_ _20038_/A VGND VGND VPWR VPWR _21932_/B sky130_fd_sc_hd__inv_2
XFILLER_101_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24915_ _24923_/CLK _24915_/D HRESETn VGND VGND VPWR VPWR _24915_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_236_0_HCLK clkbuf_8_237_0_HCLK/A VGND VGND VPWR VPWR _23744_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_46_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24051__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14929__A _24273_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12860_ _22980_/A VGND VGND VPWR VPWR _12860_/Y sky130_fd_sc_hd__inv_2
X_24846_ _24841_/CLK _24846_/D HRESETn VGND VGND VPWR VPWR _24846_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23026__B _23026_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11811_ _11803_/B VGND VGND VPWR VPWR _11811_/Y sky130_fd_sc_hd__inv_2
X_12791_ _22891_/A VGND VGND VPWR VPWR _12791_/Y sky130_fd_sc_hd__inv_2
XPHY_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24777_ _23618_/CLK _14337_/X HRESETn VGND VGND VPWR VPWR _24777_/Q sky130_fd_sc_hd__dfrtp_4
X_21989_ _21988_/X VGND VGND VPWR VPWR _21989_/Y sky130_fd_sc_hd__inv_2
XPHY_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14529_/X VGND VGND VPWR VPWR _21202_/A sky130_fd_sc_hd__buf_2
XPHY_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11741_/X VGND VGND VPWR VPWR _11743_/A sky130_fd_sc_hd__buf_2
XPHY_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23728_ _24161_/CLK _20561_/Y HRESETn VGND VGND VPWR VPWR _13526_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17194__A3 _23682_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14544_/A _14542_/A _14460_/X VGND VGND VPWR VPWR _14461_/X sky130_fd_sc_hd__a21o_4
XPHY_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11673_/A VGND VGND VPWR VPWR _11673_/Y sky130_fd_sc_hd__inv_2
XPHY_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23659_ _24643_/CLK _20734_/X HRESETn VGND VGND VPWR VPWR _23659_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _16200_/A VGND VGND VPWR VPWR _16200_/Y sky130_fd_sc_hd__inv_2
XPHY_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _22355_/A _14372_/A _22355_/A _14372_/A VGND VGND VPWR VPWR _13418_/B sky130_fd_sc_hd__a2bb2o_4
X_17180_ _20385_/A _20385_/B VGND VGND VPWR VPWR _20389_/B sky130_fd_sc_hd__or2_4
XANTENNA__21278__A2 _21553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14392_ _14387_/A _14386_/Y VGND VGND VPWR VPWR _14392_/X sky130_fd_sc_hd__and2_4
XPHY_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16131_ _11944_/X _15822_/X VGND VGND VPWR VPWR _16131_/X sky130_fd_sc_hd__or2_4
X_13343_ _24992_/Q VGND VGND VPWR VPWR _13343_/Y sky130_fd_sc_hd__inv_2
X_16062_ _16061_/Y _16059_/X _11548_/X _16059_/X VGND VGND VPWR VPWR _16062_/X sky130_fd_sc_hd__a2bb2o_4
X_13274_ _13085_/A _19365_/A VGND VGND VPWR VPWR _13275_/C sky130_fd_sc_hd__or2_4
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24892__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15013_ _24705_/Q _15013_/B VGND VGND VPWR VPWR _15013_/X sky130_fd_sc_hd__or2_4
X_12225_ _12538_/B _12222_/B _12225_/C VGND VGND VPWR VPWR _12225_/X sky130_fd_sc_hd__or3_4
XFILLER_108_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15495__A _15464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14704__A1_N _14703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24821__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19821_ _19821_/A VGND VGND VPWR VPWR _19821_/X sky130_fd_sc_hd__buf_2
X_12156_ _25130_/Q _12144_/Y _12180_/B _24549_/Q VGND VGND VPWR VPWR _12160_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_123_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24139__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_46_0_HCLK clkbuf_6_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_46_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11528__A _11527_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19752_ _19752_/A VGND VGND VPWR VPWR _21166_/B sky130_fd_sc_hd__inv_2
X_12087_ _12177_/A _12085_/Y _12185_/B _24571_/Q VGND VGND VPWR VPWR _12093_/B sky130_fd_sc_hd__a2bb2o_4
X_16964_ _16959_/X _16960_/X _16962_/X _16963_/X VGND VGND VPWR VPWR _16964_/X sky130_fd_sc_hd__or4_4
X_18703_ _18702_/Y _18697_/X _18679_/X _18697_/X VGND VGND VPWR VPWR _18703_/X sky130_fd_sc_hd__a2bb2o_4
X_15915_ _16228_/A VGND VGND VPWR VPWR _15915_/X sky130_fd_sc_hd__buf_2
X_19683_ _19682_/Y _19680_/X _19617_/X _19680_/X VGND VGND VPWR VPWR _19683_/X sky130_fd_sc_hd__a2bb2o_4
X_16895_ _16780_/Y _16784_/Y _16823_/Y _16898_/B VGND VGND VPWR VPWR _16895_/X sky130_fd_sc_hd__or4_4
XANTENNA__22121__A _21064_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18634_ _18632_/Y _18633_/Y _16556_/X _18633_/Y VGND VGND VPWR VPWR _18634_/X sky130_fd_sc_hd__a2bb2o_4
X_15846_ _15846_/A VGND VGND VPWR VPWR _15846_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13462__B _13461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18565_ _16316_/Y _23841_/Q _16316_/Y _23841_/Q VGND VGND VPWR VPWR _18565_/X sky130_fd_sc_hd__a2bb2o_4
X_12989_ _12805_/Y _12992_/B VGND VGND VPWR VPWR _12989_/Y sky130_fd_sc_hd__nand2_4
X_15777_ HWDATA[17] VGND VGND VPWR VPWR _15777_/X sky130_fd_sc_hd__buf_2
XFILLER_33_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_HCLK clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_2_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17516_ _17518_/B VGND VGND VPWR VPWR _17517_/B sky130_fd_sc_hd__inv_2
X_14728_ _24706_/Q VGND VGND VPWR VPWR _14868_/B sky130_fd_sc_hd__inv_2
X_18496_ _18434_/C _18501_/B _18449_/X VGND VGND VPWR VPWR _18496_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__23703__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14659_ _14659_/A VGND VGND VPWR VPWR _14659_/Y sky130_fd_sc_hd__inv_2
X_17447_ _17446_/X VGND VGND VPWR VPWR _17447_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17378_ _17286_/Y _17373_/B _17345_/X _17375_/B VGND VGND VPWR VPWR _17378_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16287__A1_N _14937_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19117_ _23448_/Q VGND VGND VPWR VPWR _19117_/Y sky130_fd_sc_hd__inv_2
X_16329_ _16328_/Y _16326_/X _15484_/X _16326_/X VGND VGND VPWR VPWR _16329_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24909__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19048_ _23473_/Q VGND VGND VPWR VPWR _19048_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21200__A _21393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24562__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21010_ _21010_/A _21010_/B _21010_/C VGND VGND VPWR VPWR _21010_/X sky130_fd_sc_hd__and3_4
XFILLER_82_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15671__A3 _15477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22961_ _20675_/Y _22011_/A _20541_/Y _22322_/A VGND VGND VPWR VPWR _22961_/X sky130_fd_sc_hd__o22a_4
X_24700_ _24698_/CLK _24700_/D HRESETn VGND VGND VPWR VPWR _24700_/Q sky130_fd_sc_hd__dfrtp_4
X_21912_ _21924_/A _21912_/B VGND VGND VPWR VPWR _21914_/B sky130_fd_sc_hd__or2_4
XANTENNA__22941__A2 _20910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15481__A1_N _12101_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22892_ _21972_/X _22891_/X _22634_/X _24529_/Q _21187_/X VGND VGND VPWR VPWR _22892_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_55_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16081__B1 _15777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15423__A3 _15416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21870__A _21870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24631_ _23618_/CLK _24631_/D HRESETn VGND VGND VPWR VPWR _14639_/A sky130_fd_sc_hd__dfstp_4
X_21843_ _20782_/X _21839_/X _21840_/X _21843_/D VGND VGND VPWR VPWR _21843_/X sky130_fd_sc_hd__and4_4
XFILLER_3_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_66_0_HCLK clkbuf_8_67_0_HCLK/A VGND VGND VPWR VPWR _24968_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24562_ _25123_/CLK _24562_/D HRESETn VGND VGND VPWR VPWR _24562_/Q sky130_fd_sc_hd__dfrtp_4
X_21774_ _21762_/X _21774_/B VGND VGND VPWR VPWR _21774_/X sky130_fd_sc_hd__or2_4
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23513_ _23537_/CLK _23513_/D VGND VGND VPWR VPWR _18934_/A sky130_fd_sc_hd__dfxtp_4
X_20725_ _24026_/Q _24024_/Q VGND VGND VPWR VPWR _20725_/X sky130_fd_sc_hd__and2_4
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24493_ _24307_/CLK _24493_/D HRESETn VGND VGND VPWR VPWR _24493_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14484__A _14479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23444_ _23440_/CLK _23444_/D VGND VGND VPWR VPWR _17772_/B sky130_fd_sc_hd__dfxtp_4
X_20656_ _20656_/A VGND VGND VPWR VPWR _20656_/Y sky130_fd_sc_hd__inv_2
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23375_ _25002_/CLK _23375_/D VGND VGND VPWR VPWR _13309_/B sky130_fd_sc_hd__dfxtp_4
X_20587_ _20584_/Y _20579_/Y _20590_/B VGND VGND VPWR VPWR _20587_/X sky130_fd_sc_hd__o21a_4
X_25114_ _25115_/CLK _12263_/Y HRESETn VGND VGND VPWR VPWR _12127_/A sky130_fd_sc_hd__dfrtp_4
X_22326_ _22500_/A _22326_/B VGND VGND VPWR VPWR _22331_/C sky130_fd_sc_hd__nor2_4
XANTENNA__15895__B1 _15894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14698__B2 _24124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25045_ _25034_/CLK _12751_/X HRESETn VGND VGND VPWR VPWR _12568_/A sky130_fd_sc_hd__dfrtp_4
X_22257_ _21051_/X VGND VGND VPWR VPWR _22299_/A sky130_fd_sc_hd__buf_2
XANTENNA__12732__A _12749_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21968__B1 _20918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12010_ _12054_/A _12007_/X _11981_/X _12007_/X VGND VGND VPWR VPWR _25139_/D sky130_fd_sc_hd__a2bb2o_4
X_21208_ _21201_/X _21207_/X _14488_/X VGND VGND VPWR VPWR _21208_/X sky130_fd_sc_hd__o21a_4
XFILLER_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22188_ _20866_/A VGND VGND VPWR VPWR _22188_/X sky130_fd_sc_hd__buf_2
XANTENNA__24232__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21139_ _21333_/A _19774_/Y VGND VGND VPWR VPWR _21139_/X sky130_fd_sc_hd__or2_4
XFILLER_8_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13961_ _23647_/D _13960_/X _24805_/Q _23647_/D VGND VGND VPWR VPWR _24893_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15662__A3 _15320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12912_ _12884_/X _12892_/X _12788_/Y VGND VGND VPWR VPWR _12913_/C sky130_fd_sc_hd__o21a_4
X_15700_ _12335_/Y _15698_/X _15386_/X _15698_/X VGND VGND VPWR VPWR _15700_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22932__A2 _22285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16680_ _16680_/A _16032_/A _16680_/C _16679_/X VGND VGND VPWR VPWR _16680_/X sky130_fd_sc_hd__or4_4
XFILLER_100_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13892_ _13908_/A VGND VGND VPWR VPWR _13892_/X sky130_fd_sc_hd__buf_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16072__B1 _15855_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22876__A _14714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12843_ _12880_/A _22463_/A _12880_/A _22463_/A VGND VGND VPWR VPWR _12844_/D sky130_fd_sc_hd__a2bb2o_4
X_15631_ _15630_/Y _15628_/X _15279_/X _15628_/X VGND VGND VPWR VPWR _24506_/D sky130_fd_sc_hd__a2bb2o_4
X_24829_ _24824_/CLK _14183_/X HRESETn VGND VGND VPWR VPWR _24829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22595__B _21979_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15562_ _15561_/X VGND VGND VPWR VPWR _15562_/Y sky130_fd_sc_hd__inv_2
X_18350_ _16448_/A _18425_/A _16408_/Y _23839_/Q VGND VGND VPWR VPWR _18357_/B sky130_fd_sc_hd__a2bb2o_4
X_12774_ _22308_/A VGND VGND VPWR VPWR _12774_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25091__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14513_/A VGND VGND VPWR VPWR _14513_/Y sky130_fd_sc_hd__inv_2
X_17301_ _17300_/X VGND VGND VPWR VPWR _17362_/A sky130_fd_sc_hd__buf_2
XPHY_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _11725_/A VGND VGND VPWR VPWR _11725_/X sky130_fd_sc_hd__buf_2
XANTENNA__25020__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _12121_/Y _15490_/X _11573_/X _15490_/X VGND VGND VPWR VPWR _24562_/D sky130_fd_sc_hd__a2bb2o_4
X_18281_ _18278_/A _18277_/X VGND VGND VPWR VPWR _18281_/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _24745_/Q _14444_/B VGND VGND VPWR VPWR _14445_/A sky130_fd_sc_hd__and2_4
X_17232_ _11749_/X _17230_/X _13026_/X _17231_/Y VGND VGND VPWR VPWR _17233_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22448__A1 _21570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _11657_/A _11655_/Y _13557_/A _23914_/Q VGND VGND VPWR VPWR _11656_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_70_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20459__B1 _20446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17163_ _17030_/Y _17161_/X _17162_/Y VGND VGND VPWR VPWR _17163_/X sky130_fd_sc_hd__o21a_4
XFILLER_80_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14375_ _14374_/X VGND VGND VPWR VPWR _14420_/B sky130_fd_sc_hd__inv_2
XFILLER_11_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11587_ _11587_/A VGND VGND VPWR VPWR _11587_/Y sky130_fd_sc_hd__inv_2
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16114_ _24329_/Q VGND VGND VPWR VPWR _21716_/A sky130_fd_sc_hd__inv_2
X_13326_ _13326_/A VGND VGND VPWR VPWR _21707_/B sky130_fd_sc_hd__buf_2
X_17094_ _17128_/A _17043_/B _17132_/A _17124_/B VGND VGND VPWR VPWR _17116_/B sky130_fd_sc_hd__or4_4
XANTENNA__22116__A _20753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15886__B1 _15511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16045_ _16083_/A VGND VGND VPWR VPWR _16046_/A sky130_fd_sc_hd__buf_2
X_13257_ _13057_/X _13256_/X _24998_/Q _13116_/X VGND VGND VPWR VPWR _13257_/X sky130_fd_sc_hd__o22a_4
X_12208_ _12079_/X _12219_/A _12185_/B _12219_/B VGND VGND VPWR VPWR _12209_/A sky130_fd_sc_hd__or4_4
XANTENNA__21423__A2 _22279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13188_ _13110_/A _23323_/Q VGND VGND VPWR VPWR _13189_/C sky130_fd_sc_hd__or2_4
XFILLER_83_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19804_ _19800_/X _18067_/X _13665_/A _13085_/B _19802_/X VGND VGND VPWR VPWR _23205_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24022__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12139_ _12173_/C _24560_/Q _12173_/C _24560_/Q VGND VGND VPWR VPWR _12139_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19425__A _19417_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17996_ _11655_/Y _17995_/X _17202_/X _17995_/X VGND VGND VPWR VPWR _23916_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19735_ _23230_/Q VGND VGND VPWR VPWR _22100_/B sky130_fd_sc_hd__inv_2
XFILLER_133_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16947_ _16921_/C _16921_/D VGND VGND VPWR VPWR _16952_/B sky130_fd_sc_hd__or2_4
XANTENNA__12368__A2_N _24480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14569__A _14569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23955__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19666_ _19530_/A _18031_/B _18020_/X _18039_/X VGND VGND VPWR VPWR _19667_/A sky130_fd_sc_hd__or4_4
XANTENNA__25179__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16878_ _16867_/A _16874_/B _16877_/X VGND VGND VPWR VPWR _24082_/D sky130_fd_sc_hd__and3_4
XANTENNA__20934__A1 _20931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20934__B2 _22439_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18617_ _18617_/A _18617_/B VGND VGND VPWR VPWR _18617_/X sky130_fd_sc_hd__or2_4
X_15829_ _15818_/Y _15827_/X _15828_/X _15827_/X VGND VGND VPWR VPWR _15829_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25108__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19597_ _19597_/A VGND VGND VPWR VPWR _19597_/X sky130_fd_sc_hd__buf_2
XFILLER_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12089__A _12089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18548_ _18427_/A _18523_/X _18482_/A _18546_/B VGND VGND VPWR VPWR _18548_/X sky130_fd_sc_hd__a211o_4
X_18479_ _18479_/A _18479_/B VGND VGND VPWR VPWR _18480_/C sky130_fd_sc_hd__or2_4
X_20510_ _20484_/X _20509_/Y _15352_/A _20488_/X VGND VGND VPWR VPWR _23715_/D sky130_fd_sc_hd__a2bb2o_4
X_21490_ _15463_/A VGND VGND VPWR VPWR _21490_/X sky130_fd_sc_hd__buf_2
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16008__B _15439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20441_ _20440_/X VGND VGND VPWR VPWR _20441_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24743__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23160_ _25112_/CLK _23160_/D VGND VGND VPWR VPWR _23160_/Q sky130_fd_sc_hd__dfxtp_4
X_20372_ _20372_/A _17176_/X VGND VGND VPWR VPWR _20372_/Y sky130_fd_sc_hd__nand2_4
X_22111_ _20975_/A _22109_/X _22111_/C VGND VGND VPWR VPWR _22111_/X sky130_fd_sc_hd__and3_4
X_23091_ _23939_/CLK _20104_/X VGND VGND VPWR VPWR _23091_/Q sky130_fd_sc_hd__dfxtp_4
X_22042_ _23085_/Q _22042_/B VGND VGND VPWR VPWR _22042_/X sky130_fd_sc_hd__or2_4
XANTENNA__21865__A _21864_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22611__B2 _22531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15629__B1 _15393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19549__A2_N _19546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14301__B1 _14213_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23993_ _23993_/CLK _23993_/D HRESETn VGND VGND VPWR VPWR _17310_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14479__A _14479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23696__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22944_ _12812_/Y _15578_/B _16710_/Y _22191_/X VGND VGND VPWR VPWR _22944_/X sky130_fd_sc_hd__o22a_4
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22875_ _22851_/X _22856_/X _22874_/X VGND VGND VPWR VPWR HRDATA[26] sky130_fd_sc_hd__a21o_4
X_24614_ _24185_/CLK _24614_/D HRESETn VGND VGND VPWR VPWR _24614_/Q sky130_fd_sc_hd__dfrtp_4
X_21826_ _20978_/A _21826_/B VGND VGND VPWR VPWR _21826_/X sky130_fd_sc_hd__or2_4
XFILLER_71_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24545_ _24545_/CLK _15526_/X HRESETn VGND VGND VPWR VPWR _24545_/Q sky130_fd_sc_hd__dfrtp_4
X_21757_ _21754_/Y _21755_/X _21701_/X _21756_/X VGND VGND VPWR VPWR _23034_/B sky130_fd_sc_hd__a211o_4
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11510_ _15314_/A _11951_/B VGND VGND VPWR VPWR _11514_/A sky130_fd_sc_hd__or2_4
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20708_ _23811_/Q _23809_/Q _23810_/Q _20707_/X VGND VGND VPWR VPWR _20708_/X sky130_fd_sc_hd__o22a_4
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12490_ _12460_/A _12488_/X _12490_/C VGND VGND VPWR VPWR _25085_/D sky130_fd_sc_hd__and3_4
X_24476_ _24307_/CLK _15697_/X HRESETn VGND VGND VPWR VPWR _12346_/A sky130_fd_sc_hd__dfrtp_4
X_21688_ _14494_/X _21688_/B _21687_/X VGND VGND VPWR VPWR _21688_/X sky130_fd_sc_hd__or3_4
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23427_ _25067_/CLK _23427_/D VGND VGND VPWR VPWR _19177_/A sky130_fd_sc_hd__dfxtp_4
X_20639_ _20639_/A VGND VGND VPWR VPWR _20644_/B sky130_fd_sc_hd__inv_2
XANTENNA__21102__A1 _16621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24484__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14160_ _14160_/A _14160_/B _14159_/Y _14155_/X VGND VGND VPWR VPWR _14160_/X sky130_fd_sc_hd__or4_4
X_23358_ _23350_/CLK _23358_/D VGND VGND VPWR VPWR _13028_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24413__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13111_ _11753_/A _13108_/X _13111_/C VGND VGND VPWR VPWR _13112_/C sky130_fd_sc_hd__and3_4
X_22309_ _12508_/A _22178_/X _24038_/Q _22260_/X VGND VGND VPWR VPWR _22310_/D sky130_fd_sc_hd__a2bb2o_4
X_14091_ _14079_/A VGND VGND VPWR VPWR _14091_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_111_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_223_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_23289_ _23288_/CLK _23289_/D VGND VGND VPWR VPWR _23289_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_106_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13042_ _13042_/A _23134_/Q VGND VGND VPWR VPWR _13043_/C sky130_fd_sc_hd__or2_4
XFILLER_4_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25028_ _25021_/CLK _12929_/X HRESETn VGND VGND VPWR VPWR _22769_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_117_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16869__A _16858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15773__A _15767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17850_ _17914_/A _17848_/X _17850_/C VGND VGND VPWR VPWR _17851_/C sky130_fd_sc_hd__and3_4
XFILLER_121_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16293__B1 _16216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16801_ _15841_/Y _24085_/Q _24415_/Q _16800_/Y VGND VGND VPWR VPWR _16801_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17781_ _17781_/A _23420_/Q VGND VGND VPWR VPWR _17783_/B sky130_fd_sc_hd__or2_4
XFILLER_93_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14993_ _15016_/A _14989_/B _14992_/X VGND VGND VPWR VPWR _14994_/A sky130_fd_sc_hd__or3_4
XFILLER_130_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19520_ _19520_/A VGND VGND VPWR VPWR _21517_/B sky130_fd_sc_hd__inv_2
XANTENNA__14843__B2 _24144_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16732_ _15945_/Y _23964_/Q _22239_/A _17490_/A VGND VGND VPWR VPWR _16739_/A sky130_fd_sc_hd__a2bb2o_4
X_13944_ _24891_/Q _13944_/B _24892_/Q VGND VGND VPWR VPWR _13944_/X sky130_fd_sc_hd__or3_4
XFILLER_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19451_ _19451_/A VGND VGND VPWR VPWR _21657_/B sky130_fd_sc_hd__inv_2
X_13875_ _13835_/X VGND VGND VPWR VPWR _13876_/D sky130_fd_sc_hd__inv_2
X_16663_ _16643_/A VGND VGND VPWR VPWR _16663_/X sky130_fd_sc_hd__buf_2
XANTENNA__15311__A1_N _21581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25201__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18402_ _16467_/Y _23816_/Q _16471_/A _18551_/A VGND VGND VPWR VPWR _18402_/X sky130_fd_sc_hd__a2bb2o_4
X_12826_ _21055_/A VGND VGND VPWR VPWR _12826_/Y sky130_fd_sc_hd__inv_2
X_15614_ _15611_/X _15599_/X _15497_/X _24517_/Q _15612_/X VGND VGND VPWR VPWR _24517_/D
+ sky130_fd_sc_hd__a32o_4
X_19382_ _19380_/Y _19378_/X _19381_/X _19378_/X VGND VGND VPWR VPWR _19382_/X sky130_fd_sc_hd__a2bb2o_4
X_16594_ _16594_/A VGND VGND VPWR VPWR _16594_/Y sky130_fd_sc_hd__inv_2
X_18333_ _18299_/X VGND VGND VPWR VPWR _18333_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12757_ _12737_/X VGND VGND VPWR VPWR _12758_/B sky130_fd_sc_hd__inv_2
X_15545_ _19445_/A VGND VGND VPWR VPWR _15545_/X sky130_fd_sc_hd__buf_2
XFILLER_128_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11708_/A _11708_/B VGND VGND VPWR VPWR _11708_/X sky130_fd_sc_hd__or2_4
X_15476_ _12089_/Y _15472_/X _11540_/X _15475_/X VGND VGND VPWR VPWR _24572_/D sky130_fd_sc_hd__a2bb2o_4
X_18264_ _18206_/X _18272_/B VGND VGND VPWR VPWR _18265_/B sky130_fd_sc_hd__or2_4
X_12688_ _12550_/X _12691_/B _12666_/X VGND VGND VPWR VPWR _12688_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14427_ _14424_/B _14412_/X _13608_/X _14426_/Y VGND VGND VPWR VPWR _24753_/D sky130_fd_sc_hd__o22a_4
X_17215_ _17215_/A VGND VGND VPWR VPWR _17215_/Y sky130_fd_sc_hd__inv_2
X_11639_ _11533_/X _15920_/A _13398_/A _25191_/Q _11537_/X VGND VGND VPWR VPWR _11639_/X
+ sky130_fd_sc_hd__a32o_4
X_18195_ _18459_/A VGND VGND VPWR VPWR _18262_/A sky130_fd_sc_hd__buf_2
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14358_ _13837_/X VGND VGND VPWR VPWR _14359_/C sky130_fd_sc_hd__inv_2
X_17146_ _17034_/A _17145_/X _17057_/X VGND VGND VPWR VPWR _17146_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_7_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22841__A1 _21490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22841__B2 _22840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24154__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13309_ _13309_/A _13309_/B VGND VGND VPWR VPWR _13310_/C sky130_fd_sc_hd__or2_4
X_17077_ _17077_/A _17076_/X VGND VGND VPWR VPWR _17077_/X sky130_fd_sc_hd__or2_4
X_14289_ _14286_/Y _14288_/X _14228_/X _14288_/X VGND VGND VPWR VPWR _14289_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15323__A2 _15319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16028_ _19189_/B VGND VGND VPWR VPWR _19144_/B sky130_fd_sc_hd__buf_2
XFILLER_48_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16284__B1 _15890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_16_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_33_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17979_ _17973_/X VGND VGND VPWR VPWR _17979_/X sky130_fd_sc_hd__buf_2
XFILLER_38_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19718_ _19709_/Y VGND VGND VPWR VPWR _19718_/X sky130_fd_sc_hd__buf_2
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19222__B1 _19221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20990_ _20994_/A _20990_/B VGND VGND VPWR VPWR _20990_/X sky130_fd_sc_hd__or2_4
XFILLER_81_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16036__B1 _13480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19773__B2 _19772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19649_ _23261_/Q VGND VGND VPWR VPWR _21935_/B sky130_fd_sc_hd__inv_2
XANTENNA__11608__A1_N _11606_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22660_ _22360_/X _22631_/X _22636_/X _22649_/X _22659_/X VGND VGND VPWR VPWR _22660_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_41_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24995__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21611_ _21606_/X _21610_/X _18048_/X VGND VGND VPWR VPWR _21611_/X sky130_fd_sc_hd__o21a_4
XFILLER_59_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22124__A3 _21981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21724__A1_N _13370_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22591_ _22591_/A _22757_/B VGND VGND VPWR VPWR _22591_/X sky130_fd_sc_hd__or2_4
XANTENNA__24924__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24330_ _24333_/CLK _16113_/X HRESETn VGND VGND VPWR VPWR _16111_/A sky130_fd_sc_hd__dfrtp_4
X_21542_ _21848_/B VGND VGND VPWR VPWR _21543_/A sky130_fd_sc_hd__buf_2
XFILLER_90_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_5_16_0_HCLK_A clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24261_ _24654_/CLK _16285_/X HRESETn VGND VGND VPWR VPWR _24261_/Q sky130_fd_sc_hd__dfrtp_4
X_21473_ _21339_/A _21465_/X _21472_/X VGND VGND VPWR VPWR _21473_/X sky130_fd_sc_hd__or3_4
XFILLER_119_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14762__A _24695_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23212_ _23308_/CLK _23212_/D VGND VGND VPWR VPWR _23212_/Q sky130_fd_sc_hd__dfxtp_4
X_20424_ _20424_/A VGND VGND VPWR VPWR _20424_/Y sky130_fd_sc_hd__inv_2
X_24192_ _24192_/CLK _16470_/X HRESETn VGND VGND VPWR VPWR _24192_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23143_ _25044_/CLK _19966_/X VGND VGND VPWR VPWR _23143_/Q sky130_fd_sc_hd__dfxtp_4
X_20355_ _14055_/Y _20344_/X _20401_/A _20354_/X VGND VGND VPWR VPWR _20355_/X sky130_fd_sc_hd__a211o_4
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23074_ _23993_/CLK _23074_/D VGND VGND VPWR VPWR _20140_/A sky130_fd_sc_hd__dfxtp_4
X_20286_ _13934_/A VGND VGND VPWR VPWR _20286_/X sky130_fd_sc_hd__buf_2
XFILLER_103_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21399__B2 _22548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23877__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22025_ _14223_/Y _20818_/X _14247_/A _21868_/B VGND VGND VPWR VPWR _22025_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22203__B _22163_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16275__B1 _24267_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11639__A1 _11533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11990_ _11990_/A VGND VGND VPWR VPWR _11990_/X sky130_fd_sc_hd__buf_2
X_23976_ _24962_/CLK _17471_/X HRESETn VGND VGND VPWR VPWR _23976_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20939__A _20777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22927_ _22334_/A _22924_/X _22927_/C VGND VGND VPWR VPWR _22938_/B sky130_fd_sc_hd__and3_4
XFILLER_72_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13660_ _22214_/A _13657_/X _11604_/X _13657_/X VGND VGND VPWR VPWR _24934_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12370__A1_N _12415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23034__B _23034_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22858_ _22858_/A VGND VGND VPWR VPWR _22858_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_36_0_HCLK clkbuf_6_18_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_36_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12611_ _12604_/X _12606_/X _12608_/X _12611_/D VGND VGND VPWR VPWR _12632_/B sky130_fd_sc_hd__or4_4
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21809_ _20961_/A _21809_/B VGND VGND VPWR VPWR _21810_/C sky130_fd_sc_hd__or2_4
X_13591_ _13591_/A _13559_/X VGND VGND VPWR VPWR _13591_/Y sky130_fd_sc_hd__nand2_4
XFILLER_73_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_99_0_HCLK clkbuf_7_99_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_99_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22789_ _15342_/Y _21562_/A _16495_/Y _21576_/X VGND VGND VPWR VPWR _22789_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24665__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15330_ _15329_/Y _15327_/X _11525_/X _15327_/X VGND VGND VPWR VPWR _24613_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12542_ _25048_/Q VGND VGND VPWR VPWR _12649_/C sky130_fd_sc_hd__inv_2
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24528_ _24478_/CLK _15595_/X HRESETn VGND VGND VPWR VPWR _24528_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15261_ _13728_/X _15260_/X _15256_/X _13726_/X _15254_/X VGND VGND VPWR VPWR _15261_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15768__A _15767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12473_ _12472_/X VGND VGND VPWR VPWR _12473_/Y sky130_fd_sc_hd__inv_2
X_24459_ _24459_/CLK _24459_/D HRESETn VGND VGND VPWR VPWR _24459_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16686__A1_N _24366_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14212_ _13921_/A _14199_/B VGND VGND VPWR VPWR _14212_/X sky130_fd_sc_hd__or2_4
X_17000_ _16186_/Y _24040_/Q _16186_/Y _24040_/Q VGND VGND VPWR VPWR _17000_/X sky130_fd_sc_hd__a2bb2o_4
X_15192_ _15192_/A _15192_/B _15192_/C VGND VGND VPWR VPWR _15192_/X sky130_fd_sc_hd__and3_4
XFILLER_32_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_HCLK clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_3_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_14143_ _24841_/Q _13492_/X _14127_/X _24987_/Q _14126_/A VGND VGND VPWR VPWR _24841_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_4_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14074_ _14074_/A _14067_/X _15236_/A _14074_/D VGND VGND VPWR VPWR _14074_/X sky130_fd_sc_hd__or4_4
X_18951_ _18949_/Y _18945_/X _18883_/X _18950_/X VGND VGND VPWR VPWR _23508_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13025_ _11733_/A VGND VGND VPWR VPWR _13271_/A sky130_fd_sc_hd__inv_2
X_17902_ _17934_/A _18934_/A VGND VGND VPWR VPWR _17904_/B sky130_fd_sc_hd__or2_4
XFILLER_79_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18882_ _18882_/A VGND VGND VPWR VPWR _18882_/Y sky130_fd_sc_hd__inv_2
X_17833_ _17927_/A _23531_/Q VGND VGND VPWR VPWR _17833_/X sky130_fd_sc_hd__or2_4
XFILLER_43_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11536__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23000__A1 _15463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15008__A _14703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17764_ _17689_/X _17764_/B _17763_/X VGND VGND VPWR VPWR _17764_/X sky130_fd_sc_hd__and3_4
XANTENNA__23000__B2 _15824_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14976_ _15123_/B VGND VGND VPWR VPWR _15094_/A sky130_fd_sc_hd__buf_2
X_19503_ _23312_/Q VGND VGND VPWR VPWR _21197_/B sky130_fd_sc_hd__inv_2
X_16715_ _24362_/Q _23944_/Q _15997_/Y _17615_/A VGND VGND VPWR VPWR _16716_/D sky130_fd_sc_hd__o22a_4
XFILLER_35_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13927_ _13927_/A _13927_/B _24887_/Q VGND VGND VPWR VPWR _13928_/B sky130_fd_sc_hd__or3_4
XFILLER_81_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17695_ _17676_/X _17693_/X _17695_/C VGND VGND VPWR VPWR _17695_/X sky130_fd_sc_hd__and3_4
XFILLER_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19434_ _13283_/B VGND VGND VPWR VPWR _19434_/Y sky130_fd_sc_hd__inv_2
X_16646_ _14751_/Y _16643_/X HWDATA[17] _16643_/X VGND VGND VPWR VPWR _24110_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13858_ _13858_/A VGND VGND VPWR VPWR _13897_/B sky130_fd_sc_hd__inv_2
XANTENNA__18038__B _17460_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12809_ _22651_/A VGND VGND VPWR VPWR _12809_/Y sky130_fd_sc_hd__inv_2
X_19365_ _19365_/A VGND VGND VPWR VPWR _19365_/Y sky130_fd_sc_hd__inv_2
X_16577_ _14823_/Y _16570_/X _16246_/X _16576_/X VGND VGND VPWR VPWR _16577_/X sky130_fd_sc_hd__a2bb2o_4
X_13789_ _13795_/A _13781_/X _13788_/X VGND VGND VPWR VPWR _13789_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22783__B _22505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18316_ _18316_/A _18303_/X VGND VGND VPWR VPWR _18317_/C sky130_fd_sc_hd__nand2_4
X_15528_ _15411_/X _15319_/Y _15432_/X _20740_/B _15527_/X VGND VGND VPWR VPWR _24544_/D
+ sky130_fd_sc_hd__a32o_4
X_19296_ _19283_/Y VGND VGND VPWR VPWR _19296_/X sky130_fd_sc_hd__buf_2
XANTENNA__24335__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18247_ _18258_/A _18221_/C _18198_/Y VGND VGND VPWR VPWR _18248_/C sky130_fd_sc_hd__o21a_4
XFILLER_50_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15459_ _15459_/A VGND VGND VPWR VPWR _15689_/A sky130_fd_sc_hd__inv_2
XANTENNA__16741__B2 _22979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18178_ _16068_/Y _23867_/Q _16102_/A _18213_/D VGND VGND VPWR VPWR _18178_/X sky130_fd_sc_hd__a2bb2o_4
X_17129_ _17129_/A _17129_/B _17128_/X VGND VGND VPWR VPWR _17129_/X sky130_fd_sc_hd__and3_4
XANTENNA__24807__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20140_ _20140_/A VGND VGND VPWR VPWR _20140_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23970__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20071_ _21181_/A _20067_/X _19963_/X _20067_/X VGND VGND VPWR VPWR _23103_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25194__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16302__A _16302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25123__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14807__B2 _24125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23830_ _23830_/CLK _23830_/D HRESETn VGND VGND VPWR VPWR _18503_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_26_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16272__A3 _16087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19613__A _19613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23780__D _20685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15848__A1_N _15846_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15480__A1 _15368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19746__B2 _19743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23761_ _24698_/CLK _23761_/D HRESETn VGND VGND VPWR VPWR _15295_/A sky130_fd_sc_hd__dfrtp_4
X_20973_ _20965_/A VGND VGND VPWR VPWR _20979_/A sky130_fd_sc_hd__buf_2
X_22712_ _22712_/A _22651_/B VGND VGND VPWR VPWR _22712_/X sky130_fd_sc_hd__and2_4
XFILLER_54_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23692_ _23668_/CLK _20252_/X HRESETn VGND VGND VPWR VPWR _20251_/A sky130_fd_sc_hd__dfrtp_4
X_22643_ _22642_/X VGND VGND VPWR VPWR _22643_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22574_ _14722_/A _22574_/B VGND VGND VPWR VPWR _22579_/B sky130_fd_sc_hd__or2_4
XANTENNA__24076__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24313_ _24049_/CLK _24313_/D HRESETn VGND VGND VPWR VPWR _24313_/Q sky130_fd_sc_hd__dfrtp_4
X_21525_ _21393_/A _21525_/B VGND VGND VPWR VPWR _21525_/X sky130_fd_sc_hd__or2_4
XFILLER_72_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24005__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16732__B2 _17490_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24244_ _24244_/CLK _16331_/X HRESETn VGND VGND VPWR VPWR _24244_/Q sky130_fd_sc_hd__dfrtp_4
X_21456_ _21455_/X VGND VGND VPWR VPWR _21457_/D sky130_fd_sc_hd__inv_2
X_20407_ _20404_/X _20406_/X _15250_/X VGND VGND VPWR VPWR _20407_/X sky130_fd_sc_hd__o21a_4
XFILLER_107_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24175_ _24177_/CLK _24175_/D HRESETn VGND VGND VPWR VPWR _24175_/Q sky130_fd_sc_hd__dfrtp_4
X_21387_ _21387_/A _21387_/B _21386_/X VGND VGND VPWR VPWR _21387_/X sky130_fd_sc_hd__and3_4
XFILLER_108_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16496__B1 _16251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23126_ _23661_/CLK _23126_/D VGND VGND VPWR VPWR _23126_/Q sky130_fd_sc_hd__dfxtp_4
X_20338_ _20333_/X _20337_/X _13916_/X VGND VGND VPWR VPWR _20338_/X sky130_fd_sc_hd__o21a_4
XFILLER_123_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23057_ _20735_/X VGND VGND VPWR VPWR IRQ[5] sky130_fd_sc_hd__buf_2
X_20269_ _14270_/A _20269_/B VGND VGND VPWR VPWR _20269_/X sky130_fd_sc_hd__and2_4
XFILLER_88_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16248__B1 _16246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23640__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22008_ _22008_/A _21868_/B VGND VGND VPWR VPWR _22008_/X sky130_fd_sc_hd__and2_4
XFILLER_62_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21792__A1 _11964_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12137__A2_N _24562_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17996__B1 _17202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21792__B2 _21791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14830_ _14805_/X _14811_/X _14820_/X _14829_/X VGND VGND VPWR VPWR _14830_/X sky130_fd_sc_hd__or4_4
XFILLER_29_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11973_ _25152_/Q VGND VGND VPWR VPWR _11973_/Y sky130_fd_sc_hd__inv_2
X_14761_ _14753_/X _14761_/B _14761_/C _14761_/D VGND VGND VPWR VPWR _14794_/A sky130_fd_sc_hd__or4_4
XFILLER_17_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23959_ _23949_/CLK _17567_/X HRESETn VGND VGND VPWR VPWR _16718_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22741__B1 _20750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24846__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16500_ _16497_/Y _16493_/X _15484_/X _16499_/X VGND VGND VPWR VPWR _16500_/X sky130_fd_sc_hd__a2bb2o_4
X_13712_ _13711_/X VGND VGND VPWR VPWR _13800_/A sky130_fd_sc_hd__buf_2
X_14692_ _14692_/A VGND VGND VPWR VPWR _24715_/D sky130_fd_sc_hd__inv_2
X_17480_ _22853_/A VGND VGND VPWR VPWR _17503_/A sky130_fd_sc_hd__inv_2
XFILLER_60_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16431_ _16430_/Y _16426_/X _16266_/X _16426_/X VGND VGND VPWR VPWR _16431_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13643_ _23036_/A VGND VGND VPWR VPWR _13643_/Y sky130_fd_sc_hd__inv_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19150_ _19148_/Y _19146_/X _19149_/X _19146_/X VGND VGND VPWR VPWR _19150_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13574_ _13574_/A VGND VGND VPWR VPWR _24961_/D sky130_fd_sc_hd__inv_2
X_16362_ _16361_/Y _16359_/X _16279_/X _16359_/X VGND VGND VPWR VPWR _16362_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18173__B1 _22401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18101_ _21648_/A _11767_/X _18100_/A _17226_/X VGND VGND VPWR VPWR _18101_/X sky130_fd_sc_hd__o22a_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _25075_/Q _12525_/B VGND VGND VPWR VPWR _12526_/C sky130_fd_sc_hd__or2_4
X_15313_ _12061_/B _15310_/X HADDR[3] _15300_/Y VGND VGND VPWR VPWR _24616_/D sky130_fd_sc_hd__a2bb2o_4
X_16293_ _14936_/Y _16286_/X _16216_/X _16247_/A VGND VGND VPWR VPWR _16293_/X sky130_fd_sc_hd__a2bb2o_4
X_19081_ _19081_/A VGND VGND VPWR VPWR _19081_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_123_0_HCLK clkbuf_7_61_0_HCLK/X VGND VGND VPWR VPWR _23872_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16723__B2 _21839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18032_ _18018_/X _18025_/X _19595_/A VGND VGND VPWR VPWR _18032_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_8_186_0_HCLK clkbuf_7_93_0_HCLK/X VGND VGND VPWR VPWR _25115_/CLK sky130_fd_sc_hd__clkbuf_1
X_12456_ _12399_/A VGND VGND VPWR VPWR _12456_/X sky130_fd_sc_hd__buf_2
X_15244_ _13764_/X _15240_/X _15243_/X VGND VGND VPWR VPWR _24649_/D sky130_fd_sc_hd__o21ai_4
XANTENNA__23799__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15175_ _15106_/A _15178_/B VGND VGND VPWR VPWR _15176_/C sky130_fd_sc_hd__nand2_4
X_12387_ _12387_/A _12387_/B _12383_/X _12387_/D VGND VGND VPWR VPWR _12397_/C sky130_fd_sc_hd__or4_4
XFILLER_125_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14126_ _14126_/A VGND VGND VPWR VPWR _14126_/X sky130_fd_sc_hd__buf_2
XFILLER_4_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16487__B1 _11536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23728__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21480__B1 _21930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19983_ _21389_/B _19982_/X _15556_/X _19982_/X VGND VGND VPWR VPWR _19983_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14057_ _24867_/Q VGND VGND VPWR VPWR _14057_/Y sky130_fd_sc_hd__inv_2
X_18934_ _18934_/A VGND VGND VPWR VPWR _18934_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22206__A2_N _11954_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16239__B1 _24285_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13008_ _12925_/X _13008_/B _13008_/C VGND VGND VPWR VPWR _13008_/X sky130_fd_sc_hd__and3_4
XANTENNA__21232__B1 _21231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18865_ _13227_/B VGND VGND VPWR VPWR _18865_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22778__B _11964_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17816_ _17816_/A _19155_/A VGND VGND VPWR VPWR _17818_/B sky130_fd_sc_hd__or2_4
XANTENNA__19490__A1_N _19486_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18796_ _18794_/Y _18790_/X _18795_/X _18790_/X VGND VGND VPWR VPWR _18796_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17747_ _17742_/A VGND VGND VPWR VPWR _17895_/A sky130_fd_sc_hd__buf_2
X_14959_ _14898_/Y _24281_/Q _24670_/Q _14958_/Y VGND VGND VPWR VPWR _14959_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21535__A1 _22146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24587__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17678_ _17694_/A _17678_/B VGND VGND VPWR VPWR _17679_/C sky130_fd_sc_hd__or2_4
XANTENNA__24516__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19417_ _19417_/A VGND VGND VPWR VPWR _19417_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16629_ _16632_/A VGND VGND VPWR VPWR _16629_/X sky130_fd_sc_hd__buf_2
XFILLER_62_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_2_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16962__B2 _24054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21299__B1 _13613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19348_ _19799_/A _18064_/X _18069_/X VGND VGND VPWR VPWR _19349_/A sky130_fd_sc_hd__or3_4
Xclkbuf_7_82_0_HCLK clkbuf_7_83_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_82_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19279_ _19279_/A VGND VGND VPWR VPWR _19279_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21310_ _14211_/Y _20826_/X _24810_/Q _21113_/C VGND VGND VPWR VPWR _21310_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22018__B _22018_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22290_ _22175_/A _22286_/Y _22349_/B _22289_/X VGND VGND VPWR VPWR _22291_/A sky130_fd_sc_hd__o22a_4
XANTENNA__16516__A1_N _16515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21241_ _21394_/A _21241_/B _21240_/X VGND VGND VPWR VPWR _21241_/X sky130_fd_sc_hd__and3_4
XANTENNA__21857__B _21745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21172_ _17639_/A VGND VGND VPWR VPWR _21172_/X sky130_fd_sc_hd__buf_2
XFILLER_104_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20123_ _20116_/X VGND VGND VPWR VPWR _20123_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20054_ _17999_/A VGND VGND VPWR VPWR _20054_/X sky130_fd_sc_hd__buf_2
X_24931_ _24974_/CLK _24931_/D HRESETn VGND VGND VPWR VPWR _24931_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17978__B1 _15497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22688__B _22574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24862_ _23657_/CLK _14080_/X HRESETn VGND VGND VPWR VPWR _14077_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23813_ _23762_/CLK _18560_/X HRESETn VGND VGND VPWR VPWR _23813_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24793_ _24859_/CLK _24793_/D HRESETn VGND VGND VPWR VPWR _24793_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22723__B1 _17502_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23744_ _23744_/CLK _23744_/D HRESETn VGND VGND VPWR VPWR _20635_/A sky130_fd_sc_hd__dfrtp_4
X_20956_ _17642_/Y VGND VGND VPWR VPWR _20962_/A sky130_fd_sc_hd__buf_2
XANTENNA__24257__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_5_31_0_HCLK_A clkbuf_5_30_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23675_ _23676_/CLK _20384_/Y HRESETn VGND VGND VPWR VPWR _23675_/Q sky130_fd_sc_hd__dfrtp_4
X_20887_ _23042_/B _20931_/A VGND VGND VPWR VPWR _20887_/Y sky130_fd_sc_hd__nand2_4
XPHY_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22626_ _22625_/X VGND VGND VPWR VPWR _22626_/Y sky130_fd_sc_hd__inv_2
XPHY_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21113__A _21097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22557_ _22992_/B VGND VGND VPWR VPWR _22557_/X sky130_fd_sc_hd__buf_2
X_12310_ _25095_/Q VGND VGND VPWR VPWR _12451_/A sky130_fd_sc_hd__inv_2
X_21508_ _21214_/A _21508_/B VGND VGND VPWR VPWR _21508_/X sky130_fd_sc_hd__or2_4
X_13290_ _11732_/B _18827_/A VGND VGND VPWR VPWR _13290_/X sky130_fd_sc_hd__or2_4
X_22488_ _16517_/Y _22488_/B VGND VGND VPWR VPWR _22488_/X sky130_fd_sc_hd__and2_4
X_12241_ _12094_/Y _12245_/B _12240_/Y VGND VGND VPWR VPWR _12241_/X sky130_fd_sc_hd__o21a_4
XANTENNA__23892__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24227_ _24197_/CLK _16377_/X HRESETn VGND VGND VPWR VPWR _16375_/A sky130_fd_sc_hd__dfrtp_4
X_21439_ _13374_/Y _20751_/X _11928_/Y _13333_/A VGND VGND VPWR VPWR _21439_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23821__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12172_ _12172_/A VGND VGND VPWR VPWR _12175_/A sky130_fd_sc_hd__inv_2
X_24158_ _24349_/CLK _16557_/X HRESETn VGND VGND VPWR VPWR _16555_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25045__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23109_ _23109_/CLK _20056_/X VGND VGND VPWR VPWR _22043_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__17038__A _24042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16980_ _16200_/A _24034_/Q _16200_/Y _17144_/A VGND VGND VPWR VPWR _16980_/X sky130_fd_sc_hd__o22a_4
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12470__A _12410_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24089_ _24088_/CLK _24089_/D HRESETn VGND VGND VPWR VPWR _24089_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22879__A _22879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15931_ _22910_/A VGND VGND VPWR VPWR _15931_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17293__A1_N _25218_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15781__A _16581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22962__B1 _20750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18650_ _18644_/Y VGND VGND VPWR VPWR _18650_/X sky130_fd_sc_hd__buf_2
XFILLER_7_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15862_ _15862_/A VGND VGND VPWR VPWR _15862_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17601_ _16712_/Y _17603_/B _17600_/Y VGND VGND VPWR VPWR _17601_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16641__B1 HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14813_ _24698_/Q _14812_/A _15033_/A _14812_/Y VGND VGND VPWR VPWR _14813_/X sky130_fd_sc_hd__o22a_4
XFILLER_92_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17984__A3 _11585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18581_ _18577_/X _18581_/B _18579_/X _18581_/D VGND VGND VPWR VPWR _18581_/X sky130_fd_sc_hd__or4_4
X_15793_ _12806_/Y _15791_/X _15386_/X _15791_/X VGND VGND VPWR VPWR _24436_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24680__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17532_ _17502_/B _17502_/D _17510_/B VGND VGND VPWR VPWR _17532_/X sky130_fd_sc_hd__or3_4
X_14744_ _14744_/A VGND VGND VPWR VPWR _14744_/Y sky130_fd_sc_hd__inv_2
X_11956_ _11955_/X VGND VGND VPWR VPWR _11956_/X sky130_fd_sc_hd__buf_2
XFILLER_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17463_ _17454_/X _17458_/Y _17462_/Y VGND VGND VPWR VPWR _17463_/X sky130_fd_sc_hd__a21o_4
X_11887_ _22006_/A _11886_/X VGND VGND VPWR VPWR _11887_/Y sky130_fd_sc_hd__nor2_4
X_14675_ _14655_/A _14674_/Y _24719_/Q _14655_/A VGND VGND VPWR VPWR _14675_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15747__A2 _15740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19202_ _19200_/Y _19196_/X _19201_/X _19196_/X VGND VGND VPWR VPWR _23418_/D sky130_fd_sc_hd__a2bb2o_4
X_16414_ _16426_/A VGND VGND VPWR VPWR _16414_/X sky130_fd_sc_hd__buf_2
X_13626_ _20847_/A VGND VGND VPWR VPWR _21448_/B sky130_fd_sc_hd__buf_2
X_17394_ _17310_/A _17393_/Y VGND VGND VPWR VPWR _17394_/X sky130_fd_sc_hd__or2_4
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19133_ _19132_/Y _19130_/X _19109_/X _19130_/X VGND VGND VPWR VPWR _23443_/D sky130_fd_sc_hd__a2bb2o_4
X_16345_ _16345_/A VGND VGND VPWR VPWR _16345_/Y sky130_fd_sc_hd__inv_2
X_13557_ _13557_/A _13557_/B VGND VGND VPWR VPWR _13558_/B sky130_fd_sc_hd__or2_4
XFILLER_9_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19242__A2_N _19239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23909__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12508_ _12508_/A _12508_/B VGND VGND VPWR VPWR _12508_/X sky130_fd_sc_hd__or2_4
X_19064_ _19071_/A VGND VGND VPWR VPWR _19064_/X sky130_fd_sc_hd__buf_2
X_13488_ _13390_/Y VGND VGND VPWR VPWR _13488_/X sky130_fd_sc_hd__buf_2
X_16276_ _16234_/A VGND VGND VPWR VPWR _16276_/X sky130_fd_sc_hd__buf_2
XFILLER_12_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18015_ _17999_/X _16228_/A _16558_/X _23040_/A _18007_/A VGND VGND VPWR VPWR _23905_/D
+ sky130_fd_sc_hd__a32o_4
X_12439_ _25097_/Q _12444_/B VGND VGND VPWR VPWR _12439_/X sky130_fd_sc_hd__or2_4
X_15227_ _15110_/B _15222_/X VGND VGND VPWR VPWR _15228_/B sky130_fd_sc_hd__nand2_4
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21453__B1 _12858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15158_ _15158_/A VGND VGND VPWR VPWR _15165_/A sky130_fd_sc_hd__buf_2
XANTENNA__19257__A2_N _19251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14109_ _11917_/D VGND VGND VPWR VPWR _14111_/C sky130_fd_sc_hd__inv_2
X_15089_ _14791_/X _15087_/X _15088_/Y VGND VGND VPWR VPWR _15089_/X sky130_fd_sc_hd__o21a_4
X_19966_ _19965_/Y _19960_/X _19392_/X _19960_/A VGND VGND VPWR VPWR _19966_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12380__A _24495_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18917_ _18917_/A VGND VGND VPWR VPWR _18917_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11708__B _11708_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19897_ _19897_/A VGND VGND VPWR VPWR _19897_/X sky130_fd_sc_hd__buf_2
XANTENNA__24768__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18848_ _21211_/B _18845_/X _15566_/X _18845_/X VGND VGND VPWR VPWR _23544_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18779_ _18778_/Y _18776_/X _18685_/X _18776_/X VGND VGND VPWR VPWR _18779_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20810_ _20809_/X VGND VGND VPWR VPWR _20810_/Y sky130_fd_sc_hd__inv_2
X_21790_ _14487_/X _21789_/X _14469_/X VGND VGND VPWR VPWR _21790_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24350__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20741_ _24964_/Q _20741_/B VGND VGND VPWR VPWR _20741_/X sky130_fd_sc_hd__and2_4
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23460_ _24733_/CLK _23460_/D VGND VGND VPWR VPWR _23460_/Q sky130_fd_sc_hd__dfxtp_4
X_20672_ _23755_/Q _13541_/X VGND VGND VPWR VPWR _20672_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__14780__A2_N _22857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22029__A _21544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22411_ _22407_/X _22411_/B VGND VGND VPWR VPWR _22416_/C sky130_fd_sc_hd__nor2_4
X_23391_ _23411_/CLK _19280_/X VGND VGND VPWR VPWR _19279_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_13_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23014__A1_N _12305_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25130_ _25130_/CLK _12205_/Y HRESETn VGND VGND VPWR VPWR _25130_/Q sky130_fd_sc_hd__dfrtp_4
X_22342_ _20472_/Y _20927_/X _20609_/Y _21870_/A VGND VGND VPWR VPWR _22342_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15866__A _24411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25061_ _25061_/CLK _25061_/D HRESETn VGND VGND VPWR VPWR _25061_/Q sky130_fd_sc_hd__dfrtp_4
X_22273_ _20917_/X _22271_/X _20903_/X _22272_/X VGND VGND VPWR VPWR _22274_/B sky130_fd_sc_hd__o22a_4
XFILLER_3_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_26_0_HCLK clkbuf_8_27_0_HCLK/A VGND VGND VPWR VPWR _24748_/CLK sky130_fd_sc_hd__clkbuf_1
X_24012_ _24013_/CLK _24012_/D HRESETn VGND VGND VPWR VPWR _24012_/Q sky130_fd_sc_hd__dfrtp_4
X_21224_ _21224_/A _21221_/X _21223_/X VGND VGND VPWR VPWR _21224_/X sky130_fd_sc_hd__and3_4
XFILLER_117_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_89_0_HCLK clkbuf_7_44_0_HCLK/X VGND VGND VPWR VPWR _23774_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_104_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21155_ _21155_/A _21152_/X _21154_/X VGND VGND VPWR VPWR _21155_/X sky130_fd_sc_hd__and3_4
XFILLER_8_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20106_ _21621_/B _20103_/X _19607_/A _20103_/X VGND VGND VPWR VPWR _20106_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21086_ _22014_/B VGND VGND VPWR VPWR _21720_/B sky130_fd_sc_hd__buf_2
XFILLER_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16697__A _23960_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22944__B1 _16710_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20037_ _22107_/B _20036_/X _19711_/X _20036_/X VGND VGND VPWR VPWR _20037_/X sky130_fd_sc_hd__a2bb2o_4
X_24914_ _24923_/CLK _13709_/X HRESETn VGND VGND VPWR VPWR _24914_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22211__B _15572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24438__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16623__B1 _24124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24845_ _24841_/CLK _14136_/X HRESETn VGND VGND VPWR VPWR _24845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11634__A HWDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11810_ _11809_/X VGND VGND VPWR VPWR _11823_/A sky130_fd_sc_hd__buf_2
XFILLER_2_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12790_ _22703_/A VGND VGND VPWR VPWR _12790_/Y sky130_fd_sc_hd__inv_2
X_21988_ _22155_/A _21985_/X _21986_/X _15892_/A _21987_/X VGND VGND VPWR VPWR _21988_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24091__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24776_ _24776_/CLK _14339_/X HRESETn VGND VGND VPWR VPWR _21549_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _23890_/Q VGND VGND VPWR VPWR _11741_/X sky130_fd_sc_hd__buf_2
X_20939_ _20777_/X _20939_/B VGND VGND VPWR VPWR _20939_/X sky130_fd_sc_hd__and2_4
XFILLER_96_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23727_ _24349_/CLK _20558_/Y HRESETn VGND VGND VPWR VPWR _13526_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__24020__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11670_/A _23915_/Q _13558_/A _11671_/Y VGND VGND VPWR VPWR _11682_/A sky130_fd_sc_hd__o22a_4
X_14460_ _24740_/Q _24739_/Q VGND VGND VPWR VPWR _14460_/X sky130_fd_sc_hd__and2_4
XFILLER_42_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23042__B _23042_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23658_ _24644_/CLK _20342_/X HRESETn VGND VGND VPWR VPWR _23658_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11993__A1_N _11992_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13411_ _13411_/A VGND VGND VPWR VPWR _22355_/A sky130_fd_sc_hd__inv_2
XPHY_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14391_ _24767_/Q _14390_/X _14388_/Y VGND VGND VPWR VPWR _14391_/X sky130_fd_sc_hd__o21a_4
XPHY_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22609_ _23960_/Q _22852_/A _22608_/X VGND VGND VPWR VPWR _22612_/C sky130_fd_sc_hd__a21o_4
XFILLER_35_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12465__A _12489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23589_ _23596_/CLK _18717_/X VGND VGND VPWR VPWR _23589_/Q sky130_fd_sc_hd__dfxtp_4
X_13342_ _13341_/Y _13339_/X _11616_/X _13339_/X VGND VGND VPWR VPWR _13342_/X sky130_fd_sc_hd__a2bb2o_4
X_16130_ _15411_/X _16135_/B _15912_/X _16817_/A _16129_/X VGND VGND VPWR VPWR _16130_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21778__A _21383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13273_ _13136_/A _13273_/B VGND VGND VPWR VPWR _13273_/X sky130_fd_sc_hd__or2_4
X_16061_ _16061_/A VGND VGND VPWR VPWR _16061_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15362__B1 _11573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12224_ _12184_/D _12192_/B _12171_/B VGND VGND VPWR VPWR _12225_/C sky130_fd_sc_hd__o21a_4
X_15012_ _15012_/A VGND VGND VPWR VPWR _15013_/B sky130_fd_sc_hd__inv_2
XFILLER_120_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19820_ _19820_/A VGND VGND VPWR VPWR _21781_/B sky130_fd_sc_hd__inv_2
X_12155_ _12154_/Y _24575_/Q _12154_/Y _24575_/Q VGND VGND VPWR VPWR _12160_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17654__A2 _16222_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19751_ _21349_/B _19750_/X _19728_/X _19750_/X VGND VGND VPWR VPWR _19751_/X sky130_fd_sc_hd__a2bb2o_4
X_12086_ _12086_/A VGND VGND VPWR VPWR _12185_/B sky130_fd_sc_hd__inv_2
X_16963_ _16155_/Y _17080_/A _16155_/Y _17080_/A VGND VGND VPWR VPWR _16963_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24861__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18702_ _18702_/A VGND VGND VPWR VPWR _18702_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22935__B1 _22530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15914_ _11535_/X _15410_/X _15912_/X _24393_/Q _15913_/X VGND VGND VPWR VPWR _15914_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_42_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19682_ _19682_/A VGND VGND VPWR VPWR _19682_/Y sky130_fd_sc_hd__inv_2
X_16894_ _16826_/C _16893_/X VGND VGND VPWR VPWR _16898_/B sky130_fd_sc_hd__or2_4
XANTENNA__24179__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16614__B1 _24128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18633_ _18633_/A _17222_/B VGND VGND VPWR VPWR _18633_/Y sky130_fd_sc_hd__nor2_4
X_15845_ _15844_/Y _15842_/X _11548_/X _15842_/X VGND VGND VPWR VPWR _24420_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24108__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11544__A _25216_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18564_ _16385_/Y _23814_/Q _16375_/A _18421_/B VGND VGND VPWR VPWR _18564_/X sky130_fd_sc_hd__a2bb2o_4
X_15776_ _12797_/Y _15773_/X _15775_/X _15773_/X VGND VGND VPWR VPWR _24447_/D sky130_fd_sc_hd__a2bb2o_4
X_12988_ _12992_/A _12984_/X _12987_/Y VGND VGND VPWR VPWR _12988_/X sky130_fd_sc_hd__and3_4
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20857__A _24125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17515_ _17505_/C _17515_/B _16733_/Y _17515_/D VGND VGND VPWR VPWR _17518_/B sky130_fd_sc_hd__or4_4
X_14727_ _24690_/Q _14726_/A _15067_/B _14726_/Y VGND VGND VPWR VPWR _14727_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11939_ _11939_/A VGND VGND VPWR VPWR _20847_/A sky130_fd_sc_hd__buf_2
X_18495_ _18358_/Y _18495_/B _18434_/D _18495_/D VGND VGND VPWR VPWR _18501_/B sky130_fd_sc_hd__or4_4
X_17446_ _11505_/A _20842_/B _11726_/Y _11720_/X VGND VGND VPWR VPWR _17446_/X sky130_fd_sc_hd__or4_4
X_14658_ _14612_/C _14627_/B _14612_/C _14627_/B VGND VGND VPWR VPWR _14659_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14258__A1_N _14257_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13609_ _13460_/X VGND VGND VPWR VPWR _13609_/X sky130_fd_sc_hd__buf_2
XFILLER_92_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17377_ _17390_/A _17377_/B _17376_/X VGND VGND VPWR VPWR _23999_/D sky130_fd_sc_hd__and3_4
X_14589_ _19123_/D _14589_/B VGND VGND VPWR VPWR _14589_/X sky130_fd_sc_hd__or2_4
XFILLER_14_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19116_ _19113_/Y _19114_/X _19115_/X _19114_/X VGND VGND VPWR VPWR _19116_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23743__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16328_ _24245_/Q VGND VGND VPWR VPWR _16328_/Y sky130_fd_sc_hd__inv_2
X_19047_ _19046_/Y _19042_/X _18932_/X _19042_/X VGND VGND VPWR VPWR _23474_/D sky130_fd_sc_hd__a2bb2o_4
X_16259_ HWDATA[20] VGND VGND VPWR VPWR _16259_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_242_0_HCLK clkbuf_8_243_0_HCLK/A VGND VGND VPWR VPWR _24138_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24949__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19949_ _19945_/Y _19948_/X _17993_/X _19948_/X VGND VGND VPWR VPWR _23150_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22312__A _22312_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22926__B1 _22858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13934__A _13934_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22960_ _16483_/Y _21576_/X _15329_/Y _22452_/X VGND VGND VPWR VPWR _22960_/X sky130_fd_sc_hd__o22a_4
XFILLER_110_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24531__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16605__B1 _16451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22031__B _20800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21911_ _20975_/A _21909_/X _21910_/X VGND VGND VPWR VPWR _21911_/X sky130_fd_sc_hd__and3_4
X_22891_ _22891_/A _22703_/B VGND VGND VPWR VPWR _22891_/X sky130_fd_sc_hd__or2_4
XANTENNA__22966__B _22999_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21842_ _12403_/B _22178_/A VGND VGND VPWR VPWR _21843_/D sky130_fd_sc_hd__or2_4
XFILLER_23_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24630_ _23618_/CLK _15277_/X HRESETn VGND VGND VPWR VPWR _20393_/A sky130_fd_sc_hd__dfstp_4
XFILLER_58_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14092__B1 _13638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20767__A _20931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24561_ _24545_/CLK _24561_/D HRESETn VGND VGND VPWR VPWR _24561_/Q sky130_fd_sc_hd__dfrtp_4
X_21773_ _21777_/A _18649_/Y VGND VGND VPWR VPWR _21773_/X sky130_fd_sc_hd__or2_4
XFILLER_36_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20724_ _20723_/A _20723_/B _24022_/Q _20723_/X VGND VGND VPWR VPWR _20724_/X sky130_fd_sc_hd__o22a_4
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23512_ _23537_/CLK _23512_/D VGND VGND VPWR VPWR _23512_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24492_ _24042_/CLK _15673_/X HRESETn VGND VGND VPWR VPWR _24492_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22982__A _22982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22037__A2_N _22246_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23443_ _23440_/CLK _23443_/D VGND VGND VPWR VPWR _17808_/B sky130_fd_sc_hd__dfxtp_4
X_20655_ _20647_/X _20654_/Y _24180_/Q _20651_/X VGND VGND VPWR VPWR _23749_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15592__B1 _15332_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_52_0_HCLK clkbuf_6_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_52_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23374_ _23374_/CLK _19330_/X VGND VGND VPWR VPWR _13013_/B sky130_fd_sc_hd__dfxtp_4
X_20586_ _20585_/X VGND VGND VPWR VPWR _20590_/B sky130_fd_sc_hd__buf_2
XFILLER_136_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22325_ _22322_/X _22323_/X _22280_/X _22324_/X VGND VGND VPWR VPWR _22326_/B sky130_fd_sc_hd__o22a_4
XANTENNA__15596__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25113_ _25115_/CLK _12274_/X HRESETn VGND VGND VPWR VPWR _12071_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22209__A2 _22208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19702__A2_N _19701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21417__B1 _21062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25044_ _25044_/CLK _25044_/D HRESETn VGND VGND VPWR VPWR _25044_/Q sky130_fd_sc_hd__dfrtp_4
X_22256_ _22256_/A _22256_/B VGND VGND VPWR VPWR _22256_/X sky130_fd_sc_hd__and2_4
XANTENNA__21968__A1 _20940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21207_ _21372_/A _21207_/B _21207_/C VGND VGND VPWR VPWR _21207_/X sky130_fd_sc_hd__and3_4
XANTENNA__21968__B2 _21967_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11629__A HWDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22187_ _22187_/A _22153_/B VGND VGND VPWR VPWR _22187_/X sky130_fd_sc_hd__or2_4
XFILLER_117_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24619__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21138_ _21153_/A VGND VGND VPWR VPWR _21333_/A sky130_fd_sc_hd__buf_2
XFILLER_120_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_5_0_HCLK_A clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16962__A1_N _16202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22917__B1 _24573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13960_ _13939_/A _13944_/X _13939_/Y _13945_/Y VGND VGND VPWR VPWR _13960_/X sky130_fd_sc_hd__o22a_4
X_21069_ _21069_/A VGND VGND VPWR VPWR _21069_/X sky130_fd_sc_hd__buf_2
XANTENNA__24272__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12911_ _12911_/A VGND VGND VPWR VPWR _12922_/A sky130_fd_sc_hd__buf_2
XFILLER_47_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13891_ _13891_/A VGND VGND VPWR VPWR _13908_/A sky130_fd_sc_hd__buf_2
XANTENNA__24201__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22876__B _22745_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15630_ _15630_/A VGND VGND VPWR VPWR _15630_/Y sky130_fd_sc_hd__inv_2
X_12842_ _22474_/A VGND VGND VPWR VPWR _12880_/A sky130_fd_sc_hd__inv_2
XFILLER_73_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24828_ _24824_/CLK _14185_/X HRESETn VGND VGND VPWR VPWR _24828_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23053__A _23040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15561_ _19835_/A VGND VGND VPWR VPWR _15561_/X sky130_fd_sc_hd__buf_2
X_12773_ _12773_/A VGND VGND VPWR VPWR _12773_/Y sky130_fd_sc_hd__inv_2
XPHY_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24759_ _24968_/CLK _14413_/X HRESETn VGND VGND VPWR VPWR _13413_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17505_/C VGND VGND VPWR VPWR _17300_/X sky130_fd_sc_hd__buf_2
XPHY_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _21756_/A _14480_/X _14511_/A _14484_/X VGND VGND VPWR VPWR _14513_/A sky130_fd_sc_hd__o22a_4
XANTENNA__17051__A _24058_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11724_ _14013_/A _11723_/X VGND VGND VPWR VPWR _11725_/A sky130_fd_sc_hd__and2_4
X_18280_ _18284_/A _18280_/B _18279_/Y VGND VGND VPWR VPWR _23863_/D sky130_fd_sc_hd__and3_4
XPHY_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _12117_/Y _15490_/X _11570_/X _15490_/X VGND VGND VPWR VPWR _24563_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17230_/X VGND VGND VPWR VPWR _17231_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _21871_/A VGND VGND VPWR VPWR _11655_/Y sky130_fd_sc_hd__inv_2
X_14443_ _14528_/A _14443_/B VGND VGND VPWR VPWR _14444_/B sky130_fd_sc_hd__and2_4
XPHY_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17162_ _17030_/Y _17161_/X _17057_/X VGND VGND VPWR VPWR _17162_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_127_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22177__A1_N _11606_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11586_ _11583_/Y _11577_/X _11585_/X _11577_/X VGND VGND VPWR VPWR _25204_/D sky130_fd_sc_hd__a2bb2o_4
X_14374_ _14374_/A _14373_/Y VGND VGND VPWR VPWR _14374_/X sky130_fd_sc_hd__or2_4
XANTENNA__25060__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16113_ _21858_/A _16112_/X _15894_/X _16112_/X VGND VGND VPWR VPWR _16113_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13325_ _13324_/X VGND VGND VPWR VPWR _13326_/A sky130_fd_sc_hd__buf_2
XFILLER_127_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17093_ _17093_/A VGND VGND VPWR VPWR _17093_/Y sky130_fd_sc_hd__inv_2
X_16044_ _16043_/X VGND VGND VPWR VPWR _16083_/A sky130_fd_sc_hd__buf_2
XANTENNA__21020__B _21020_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13256_ _11710_/X _13240_/X _13255_/X _24999_/Q _13114_/X VGND VGND VPWR VPWR _13256_/X
+ sky130_fd_sc_hd__o32a_4
X_12207_ _12207_/A _12207_/B VGND VGND VPWR VPWR _12219_/B sky130_fd_sc_hd__or2_4
X_13187_ _13219_/A _13187_/B VGND VGND VPWR VPWR _13189_/B sky130_fd_sc_hd__or2_4
XFILLER_9_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_72_0_HCLK clkbuf_7_36_0_HCLK/X VGND VGND VPWR VPWR _24974_/CLK sky130_fd_sc_hd__clkbuf_1
X_12138_ _25117_/Q VGND VGND VPWR VPWR _12173_/C sky130_fd_sc_hd__inv_2
X_19803_ _19800_/X _18067_/X _13663_/A _23206_/Q _19802_/X VGND VGND VPWR VPWR _19803_/X
+ sky130_fd_sc_hd__a32o_4
X_17995_ _17975_/Y VGND VGND VPWR VPWR _17995_/X sky130_fd_sc_hd__buf_2
XANTENNA__22908__B1 _24423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12069_ _12069_/A VGND VGND VPWR VPWR _20889_/A sky130_fd_sc_hd__inv_2
X_16946_ _16946_/A VGND VGND VPWR VPWR _16946_/Y sky130_fd_sc_hd__inv_2
X_19734_ _19733_/Y _19727_/X _19641_/X _19709_/Y VGND VGND VPWR VPWR _23231_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21971__A _20814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19665_ _19665_/A VGND VGND VPWR VPWR _22085_/B sky130_fd_sc_hd__inv_2
X_16877_ _16821_/A _16881_/B VGND VGND VPWR VPWR _16877_/X sky130_fd_sc_hd__or2_4
XFILLER_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18616_ _18616_/A _18616_/B VGND VGND VPWR VPWR _18617_/B sky130_fd_sc_hd__or2_4
X_15828_ HWDATA[31] VGND VGND VPWR VPWR _15828_/X sky130_fd_sc_hd__buf_2
XFILLER_53_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19596_ _19613_/A VGND VGND VPWR VPWR _19596_/X sky130_fd_sc_hd__buf_2
XANTENNA__23995__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18547_ _18540_/A _18543_/B _18547_/C VGND VGND VPWR VPWR _23818_/D sky130_fd_sc_hd__and3_4
X_15759_ _15748_/X _15740_/X _15477_/X _24455_/Q _15746_/X VGND VGND VPWR VPWR _24455_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23924__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18478_ _18468_/X VGND VGND VPWR VPWR _18479_/B sky130_fd_sc_hd__inv_2
XANTENNA__25148__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17429_ _17429_/A VGND VGND VPWR VPWR _17430_/B sky130_fd_sc_hd__inv_2
XFILLER_53_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20440_ _21728_/A _20437_/X _20425_/X _20439_/X VGND VGND VPWR VPWR _20440_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22307__A _22307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20371_ _20371_/A VGND VGND VPWR VPWR _20371_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16669__A3 _15704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16305__A _16305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22110_ _20966_/A _22110_/B VGND VGND VPWR VPWR _22111_/C sky130_fd_sc_hd__or2_4
XFILLER_106_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23090_ _23939_/CLK _20106_/X VGND VGND VPWR VPWR _20105_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_115_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24783__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22041_ _21582_/X VGND VGND VPWR VPWR _22041_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24712__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16146__A2_N _16138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23992_ _23992_/CLK _23992_/D HRESETn VGND VGND VPWR VPWR _17311_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_99_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22914__A3 _22459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22943_ _22943_/A _22942_/X VGND VGND VPWR VPWR _22943_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__19240__B2 _19239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22696__B _22587_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14065__B1 _13645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22127__A1 _22155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22874_ _22997_/A _22874_/B _22874_/C _22873_/Y VGND VGND VPWR VPWR _22874_/X sky130_fd_sc_hd__or4_4
X_24613_ _24612_/CLK _24613_/D HRESETn VGND VGND VPWR VPWR _15329_/A sky130_fd_sc_hd__dfrtp_4
X_21825_ _20975_/A _21825_/B _21824_/X VGND VGND VPWR VPWR _21825_/X sky130_fd_sc_hd__and3_4
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21756_ _21756_/A _21756_/B VGND VGND VPWR VPWR _21756_/X sky130_fd_sc_hd__and2_4
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24544_ _24017_/CLK _24544_/D HRESETn VGND VGND VPWR VPWR _20740_/B sky130_fd_sc_hd__dfrtp_4
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20707_ _23811_/Q _23809_/Q VGND VGND VPWR VPWR _20707_/X sky130_fd_sc_hd__and2_4
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21687_ _21682_/X _21686_/X _14440_/X VGND VGND VPWR VPWR _21687_/X sky130_fd_sc_hd__o21a_4
XFILLER_138_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24475_ _24307_/CLK _15699_/X HRESETn VGND VGND VPWR VPWR _12329_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20638_ _13537_/C _13524_/D VGND VGND VPWR VPWR _20639_/A sky130_fd_sc_hd__or2_4
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23426_ _25067_/CLK _19180_/X VGND VGND VPWR VPWR _23426_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22217__A _11529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23357_ _23350_/CLK _23357_/D VGND VGND VPWR VPWR _13104_/B sky130_fd_sc_hd__dfxtp_4
X_20569_ _20568_/X VGND VGND VPWR VPWR _23730_/D sky130_fd_sc_hd__inv_2
XFILLER_50_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13110_ _13110_/A _19470_/A VGND VGND VPWR VPWR _13111_/C sky130_fd_sc_hd__or2_4
X_22308_ _22308_/A _22299_/A VGND VGND VPWR VPWR _22308_/X sky130_fd_sc_hd__and2_4
XFILLER_125_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14090_ _14090_/A VGND VGND VPWR VPWR _14090_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16729__A2_N _16718_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23288_ _23288_/CLK _23288_/D VGND VGND VPWR VPWR _23288_/Q sky130_fd_sc_hd__dfxtp_4
X_13041_ _13045_/A _13041_/B VGND VGND VPWR VPWR _13043_/B sky130_fd_sc_hd__or2_4
X_22239_ _22239_/A _22238_/X VGND VGND VPWR VPWR _22239_/X sky130_fd_sc_hd__or2_4
XFILLER_3_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25027_ _24451_/CLK _12932_/Y HRESETn VGND VGND VPWR VPWR _12845_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24453__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_59_0_HCLK clkbuf_7_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_59_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16800_ _24079_/Q VGND VGND VPWR VPWR _16800_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17780_ _17780_/A _17778_/X _17780_/C VGND VGND VPWR VPWR _17784_/B sky130_fd_sc_hd__and3_4
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20548__A1_N _20419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14992_ _14881_/X _14982_/X _14882_/A VGND VGND VPWR VPWR _14992_/X sky130_fd_sc_hd__o21a_4
XFILLER_130_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16731_ _16731_/A _16728_/X _16729_/X _16730_/X VGND VGND VPWR VPWR _16731_/X sky130_fd_sc_hd__or4_4
XFILLER_75_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13943_ _13928_/C _13943_/B _24890_/Q VGND VGND VPWR VPWR _13944_/B sky130_fd_sc_hd__or3_4
X_19450_ _19447_/Y _19441_/X _19448_/X _19449_/X VGND VGND VPWR VPWR _23332_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16662_ _14744_/Y _16659_/X _16451_/X _16659_/X VGND VGND VPWR VPWR _16662_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13874_ _13828_/C VGND VGND VPWR VPWR _13880_/B sky130_fd_sc_hd__inv_2
XANTENNA__14056__B1 _13632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18401_ _18394_/X _18401_/B _18401_/C _18401_/D VGND VGND VPWR VPWR _18401_/X sky130_fd_sc_hd__or4_4
X_15613_ _15611_/X _15599_/X _15494_/X _24518_/Q _15612_/X VGND VGND VPWR VPWR _24518_/D
+ sky130_fd_sc_hd__a32o_4
X_12825_ _12951_/A _12823_/Y _21840_/A _21851_/A VGND VGND VPWR VPWR _12825_/X sky130_fd_sc_hd__a2bb2o_4
X_19381_ _11625_/A VGND VGND VPWR VPWR _19381_/X sky130_fd_sc_hd__buf_2
X_16593_ _14812_/Y _16587_/X _16179_/X _16587_/X VGND VGND VPWR VPWR _24141_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12606__B2 _24525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18332_ _18327_/X _18332_/B _18319_/X VGND VGND VPWR VPWR _23847_/D sky130_fd_sc_hd__and3_4
XFILLER_76_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15544_ _19448_/A VGND VGND VPWR VPWR _15544_/Y sky130_fd_sc_hd__inv_2
X_12756_ _12739_/X _12754_/Y _12755_/X VGND VGND VPWR VPWR _12756_/X sky130_fd_sc_hd__and3_4
XPHY_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11707_/A VGND VGND VPWR VPWR _11708_/A sky130_fd_sc_hd__buf_2
X_18263_ _18263_/A _18263_/B VGND VGND VPWR VPWR _18272_/B sky130_fd_sc_hd__or2_4
XFILLER_128_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ _15472_/A VGND VGND VPWR VPWR _15475_/X sky130_fd_sc_hd__buf_2
X_12687_ _12571_/Y _12694_/B VGND VGND VPWR VPWR _12691_/B sky130_fd_sc_hd__or2_4
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17214_ _17212_/Y _17213_/X _16671_/X _17213_/X VGND VGND VPWR VPWR _24014_/D sky130_fd_sc_hd__a2bb2o_4
X_14426_ _14424_/B VGND VGND VPWR VPWR _14426_/Y sky130_fd_sc_hd__inv_2
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11638_ HWDATA[1] VGND VGND VPWR VPWR _13398_/A sky130_fd_sc_hd__buf_2
X_18194_ _18468_/C VGND VGND VPWR VPWR _18459_/A sky130_fd_sc_hd__buf_2
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17145_ _17145_/A _17145_/B VGND VGND VPWR VPWR _17145_/X sky130_fd_sc_hd__or2_4
X_14357_ _13833_/X _14357_/B _14357_/C VGND VGND VPWR VPWR _14361_/C sky130_fd_sc_hd__or3_4
XFILLER_129_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11569_ _11541_/X VGND VGND VPWR VPWR _11569_/X sky130_fd_sc_hd__buf_2
XFILLER_128_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13308_ _13182_/A _13308_/B VGND VGND VPWR VPWR _13308_/X sky130_fd_sc_hd__or2_4
X_17076_ _17076_/A _17044_/X _17053_/A VGND VGND VPWR VPWR _17076_/X sky130_fd_sc_hd__or3_4
XFILLER_116_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14288_ _14288_/A VGND VGND VPWR VPWR _14288_/X sky130_fd_sc_hd__buf_2
XFILLER_109_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15323__A3 _15320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16027_ _16027_/A _16680_/A VGND VGND VPWR VPWR _16027_/X sky130_fd_sc_hd__or2_4
XFILLER_115_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13239_ _13207_/A _13239_/B _13239_/C VGND VGND VPWR VPWR _13240_/C sky130_fd_sc_hd__or3_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24194__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24123__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17978_ _22484_/A _17977_/X _15497_/X _17977_/X VGND VGND VPWR VPWR _23925_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16929_ _16834_/C _16932_/B _16849_/X VGND VGND VPWR VPWR _16929_/Y sky130_fd_sc_hd__a21oi_4
X_19717_ _11837_/A VGND VGND VPWR VPWR _19717_/X sky130_fd_sc_hd__buf_2
XFILLER_65_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16036__A1 _21257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19648_ _22110_/B _19647_/X _19597_/X _19647_/X VGND VGND VPWR VPWR _19648_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19579_ _19578_/Y _19576_/X _19445_/X _19576_/X VGND VGND VPWR VPWR _23285_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16807__A1_N _24423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21610_ _17644_/A _21610_/B _21609_/X VGND VGND VPWR VPWR _21610_/X sky130_fd_sc_hd__and3_4
XFILLER_0_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22590_ _22348_/X _22580_/X _22583_/X _22585_/X _22589_/Y VGND VGND VPWR VPWR _22614_/B
+ sky130_fd_sc_hd__a32o_4
X_21541_ _13614_/X VGND VGND VPWR VPWR _21848_/B sky130_fd_sc_hd__buf_2
XFILLER_90_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24260_ _24654_/CLK _16287_/X HRESETn VGND VGND VPWR VPWR _24260_/Q sky130_fd_sc_hd__dfrtp_4
X_21472_ _21468_/X _21471_/X _17639_/X VGND VGND VPWR VPWR _21472_/X sky130_fd_sc_hd__o21a_4
XFILLER_53_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24964__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23211_ _23308_/CLK _23211_/D VGND VGND VPWR VPWR _23211_/Q sky130_fd_sc_hd__dfxtp_4
X_20423_ _15403_/Y _20416_/X _20419_/X _20422_/Y VGND VGND VPWR VPWR _20424_/A sky130_fd_sc_hd__o22a_4
XANTENNA__22293__B1 _22270_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24191_ _24222_/CLK _16472_/X HRESETn VGND VGND VPWR VPWR _16471_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_119_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23142_ _23332_/CLK _19971_/X VGND VGND VPWR VPWR _23142_/Q sky130_fd_sc_hd__dfxtp_4
X_20354_ _17174_/B _20353_/Y _20349_/X VGND VGND VPWR VPWR _20354_/X sky130_fd_sc_hd__and3_4
XFILLER_122_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23073_ _23993_/CLK _20144_/X VGND VGND VPWR VPWR _23073_/Q sky130_fd_sc_hd__dfxtp_4
X_20285_ _20285_/A VGND VGND VPWR VPWR _23631_/D sky130_fd_sc_hd__inv_2
XANTENNA__21595__B _20931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22024_ _20195_/A _22024_/B VGND VGND VPWR VPWR _22028_/A sky130_fd_sc_hd__and2_4
XFILLER_0_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23975_ _23898_/CLK _23975_/D HRESETn VGND VGND VPWR VPWR _21799_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_99_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23846__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22926_ _24153_/Q _15919_/X _22858_/X _22925_/X VGND VGND VPWR VPWR _22927_/C sky130_fd_sc_hd__a211o_4
XANTENNA__14038__B1 _13638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17313__B _17270_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15786__B1 _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22857_ _22857_/A _22857_/B VGND VGND VPWR VPWR _22862_/B sky130_fd_sc_hd__or2_4
X_12610_ _12609_/Y _24517_/Q _12609_/Y _24517_/Q VGND VGND VPWR VPWR _12611_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11642__A _13644_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21808_ _22087_/A _21808_/B VGND VGND VPWR VPWR _21808_/X sky130_fd_sc_hd__or2_4
XFILLER_31_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ _13562_/B _13580_/X _13589_/Y _13587_/X _11679_/A VGND VGND VPWR VPWR _24955_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_71_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20126__A3 _19808_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22788_ _20524_/A _22170_/X _23751_/Q _21069_/X VGND VGND VPWR VPWR _22788_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_101_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12541_ _12540_/Y _12434_/A _24499_/Q VGND VGND VPWR VPWR _25069_/D sky130_fd_sc_hd__a21oi_4
XFILLER_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15538__B1 RsRx_S0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24527_ _24483_/CLK _15597_/X HRESETn VGND VGND VPWR VPWR _24527_/Q sky130_fd_sc_hd__dfrtp_4
X_21739_ _14206_/A _21082_/B VGND VGND VPWR VPWR _21739_/X sky130_fd_sc_hd__and2_4
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15260_ _15260_/A VGND VGND VPWR VPWR _15260_/X sky130_fd_sc_hd__buf_2
XFILLER_40_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12472_ _12385_/Y _12467_/B _12453_/X _12469_/B VGND VGND VPWR VPWR _12472_/X sky130_fd_sc_hd__a211o_4
X_24458_ _24502_/CLK _24458_/D HRESETn VGND VGND VPWR VPWR _12813_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14210__B1 _14209_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16750__A2 _16748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14211_ _14211_/A VGND VGND VPWR VPWR _14211_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21087__B2 _21720_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_22_0_HCLK clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_23409_ _23979_/CLK _19228_/X VGND VGND VPWR VPWR _19225_/A sky130_fd_sc_hd__dfxtp_4
X_15191_ _15191_/A _15191_/B VGND VGND VPWR VPWR _15192_/C sky130_fd_sc_hd__or2_4
XFILLER_137_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24389_ _24361_/CLK _24389_/D HRESETn VGND VGND VPWR VPWR _24389_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24634__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12772__B1 _12674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14142_ _14126_/A _14141_/X _13353_/A _13492_/X VGND VGND VPWR VPWR _24842_/D sky130_fd_sc_hd__o22a_4
XFILLER_125_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14073_ _13779_/X _14073_/B _13786_/Y VGND VGND VPWR VPWR _14074_/D sky130_fd_sc_hd__or3_4
X_18950_ _18958_/A VGND VGND VPWR VPWR _18950_/X sky130_fd_sc_hd__buf_2
XANTENNA__15710__B1 _15709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13024_ _13047_/A _13022_/X _13024_/C VGND VGND VPWR VPWR _13024_/X sky130_fd_sc_hd__and3_4
X_17901_ _17716_/X _17899_/X _17901_/C VGND VGND VPWR VPWR _17905_/B sky130_fd_sc_hd__and3_4
XFILLER_117_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18881_ _18879_/Y _18877_/X _18880_/X _18877_/X VGND VGND VPWR VPWR _18881_/X sky130_fd_sc_hd__a2bb2o_4
X_17832_ _17725_/A VGND VGND VPWR VPWR _17969_/A sky130_fd_sc_hd__buf_2
XFILLER_0_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22339__A1 _24267_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17763_ _16678_/X _17758_/X _17762_/X VGND VGND VPWR VPWR _17763_/X sky130_fd_sc_hd__or3_4
X_14975_ _14974_/X VGND VGND VPWR VPWR _15123_/B sky130_fd_sc_hd__buf_2
XFILLER_48_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_146_0_HCLK clkbuf_7_73_0_HCLK/X VGND VGND VPWR VPWR _23596_/CLK sky130_fd_sc_hd__clkbuf_1
X_16714_ _23944_/Q VGND VGND VPWR VPWR _17615_/A sky130_fd_sc_hd__inv_2
X_19502_ _19500_/Y _19501_/X _19459_/X _19501_/X VGND VGND VPWR VPWR _19502_/X sky130_fd_sc_hd__a2bb2o_4
X_13926_ _24884_/Q _13926_/B _13926_/C VGND VGND VPWR VPWR _13927_/B sky130_fd_sc_hd__or3_4
X_17694_ _17694_/A _23150_/Q VGND VGND VPWR VPWR _17695_/C sky130_fd_sc_hd__or2_4
XANTENNA__14029__B1 _13663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19433_ _19431_/Y _19432_/X _19387_/X _19432_/X VGND VGND VPWR VPWR _23337_/D sky130_fd_sc_hd__a2bb2o_4
X_16645_ _14722_/Y _16643_/X _16264_/X _16643_/X VGND VGND VPWR VPWR _16645_/X sky130_fd_sc_hd__a2bb2o_4
X_13857_ _13855_/Y _13856_/X _13831_/C _13830_/X VGND VGND VPWR VPWR _13858_/A sky130_fd_sc_hd__or4_4
XFILLER_50_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15024__A _14712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11552__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12808_ _12808_/A _12801_/X _12808_/C _12807_/X VGND VGND VPWR VPWR _12808_/X sky130_fd_sc_hd__or4_4
X_19364_ _19362_/Y _19363_/X _19227_/X _19363_/X VGND VGND VPWR VPWR _23361_/D sky130_fd_sc_hd__a2bb2o_4
X_16576_ _16584_/A VGND VGND VPWR VPWR _16576_/X sky130_fd_sc_hd__buf_2
X_13788_ _13787_/A _13786_/Y _13787_/Y _13786_/A VGND VGND VPWR VPWR _13788_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18715__B1 _17199_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18315_ _18290_/X _18312_/B _18314_/Y VGND VGND VPWR VPWR _18315_/X sky130_fd_sc_hd__and3_4
X_15527_ _15418_/A _15531_/B VGND VGND VPWR VPWR _15527_/X sky130_fd_sc_hd__or2_4
XFILLER_31_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12739_ _12739_/A _12739_/B VGND VGND VPWR VPWR _12739_/X sky130_fd_sc_hd__or2_4
X_19295_ _19295_/A VGND VGND VPWR VPWR _21352_/B sky130_fd_sc_hd__inv_2
XANTENNA__20522__B1 _20446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18246_ _18226_/A _18246_/B _18246_/C VGND VGND VPWR VPWR _23872_/D sky130_fd_sc_hd__and3_4
X_15458_ _15659_/B VGND VGND VPWR VPWR _15459_/A sky130_fd_sc_hd__buf_2
XFILLER_15_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_5_8_0_HCLK_A clkbuf_4_4_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14409_ _13435_/Y _14380_/X VGND VGND VPWR VPWR _14409_/Y sky130_fd_sc_hd__nand2_4
X_18177_ _18177_/A _18177_/B _18175_/X _18177_/D VGND VGND VPWR VPWR _18191_/B sky130_fd_sc_hd__or4_4
XFILLER_106_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15389_ _24590_/Q VGND VGND VPWR VPWR _21888_/A sky130_fd_sc_hd__inv_2
XANTENNA__19140__B1 _19095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24375__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17128_ _17128_/A _17126_/A VGND VGND VPWR VPWR _17128_/X sky130_fd_sc_hd__or2_4
XFILLER_89_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24304__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22027__B1 _23617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17059_ _17058_/X VGND VGND VPWR VPWR _24057_/D sky130_fd_sc_hd__inv_2
XFILLER_132_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15701__B1 _15390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20070_ _20070_/A VGND VGND VPWR VPWR _21181_/A sky130_fd_sc_hd__buf_2
XFILLER_135_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16302__B _16306_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_42_0_HCLK clkbuf_7_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_85_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15480__A2 _15461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20972_ _20972_/A _20972_/B VGND VGND VPWR VPWR _20975_/B sky130_fd_sc_hd__or2_4
X_23760_ _24698_/CLK _20155_/X HRESETn VGND VGND VPWR VPWR _15294_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_53_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25163__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22750__A1 _24347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18954__B1 _18953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22711_ _22637_/X _22708_/Y _22601_/X _22710_/X VGND VGND VPWR VPWR _22711_/X sky130_fd_sc_hd__a2bb2o_4
X_23691_ _23668_/CLK _20186_/X HRESETn VGND VGND VPWR VPWR _23691_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15232__A2 _15123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22642_ _22369_/X _22639_/X _22640_/X _11565_/A _22641_/X VGND VGND VPWR VPWR _22642_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_90_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15783__A3 _15499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22573_ _22542_/Y _22546_/Y _22573_/C _22572_/X VGND VGND VPWR VPWR HRDATA[17] sky130_fd_sc_hd__or4_4
XFILLER_22_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24312_ _24049_/CLK _24312_/D HRESETn VGND VGND VPWR VPWR _16160_/A sky130_fd_sc_hd__dfrtp_4
X_21524_ _21367_/A _21524_/B VGND VGND VPWR VPWR _21524_/X sky130_fd_sc_hd__or2_4
XANTENNA__22990__A _23023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21455_ _21079_/X _21452_/Y _11961_/X _21454_/X VGND VGND VPWR VPWR _21455_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22266__B1 _14831_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24243_ _24098_/CLK _24243_/D HRESETn VGND VGND VPWR VPWR _24243_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19131__B1 _19041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20406_ _20402_/A _20200_/Y _20202_/Y _20200_/A _20405_/X VGND VGND VPWR VPWR _20406_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20816__A1 _12322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24174_ _24177_/CLK _24174_/D HRESETn VGND VGND VPWR VPWR _24174_/Q sky130_fd_sc_hd__dfrtp_4
X_21386_ _21229_/A _19917_/Y VGND VGND VPWR VPWR _21386_/X sky130_fd_sc_hd__or2_4
XANTENNA__24045__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20337_ _20331_/A _20334_/Y _20335_/Y _14309_/X _20336_/X VGND VGND VPWR VPWR _20337_/X
+ sky130_fd_sc_hd__a32o_4
X_23125_ _23100_/CLK _20016_/X VGND VGND VPWR VPWR _20012_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22214__B _21357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22569__B2 _22322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23056_ _20717_/X VGND VGND VPWR VPWR IRQ[4] sky130_fd_sc_hd__buf_2
X_20268_ _20163_/C _20171_/B _20236_/X VGND VGND VPWR VPWR _23775_/D sky130_fd_sc_hd__a21o_4
XFILLER_7_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22007_ _25145_/Q _21881_/Y _22005_/X _22006_/Y VGND VGND VPWR VPWR _22007_/X sky130_fd_sc_hd__a211o_4
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20199_ _20179_/B _20198_/X _20185_/A _20161_/X VGND VGND VPWR VPWR _23774_/D sky130_fd_sc_hd__a211o_4
XFILLER_130_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21792__A2 _21749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22230__A _22230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14948__A _24667_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23680__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_219_0_HCLK clkbuf_8_219_0_HCLK/A VGND VGND VPWR VPWR _24098_/CLK sky130_fd_sc_hd__clkbuf_1
X_14760_ _14759_/Y _24107_/Q _14759_/Y _24107_/Q VGND VGND VPWR VPWR _14761_/D sky130_fd_sc_hd__a2bb2o_4
X_11972_ _11970_/Y _11966_/X _11620_/X _11971_/X VGND VGND VPWR VPWR _11972_/X sky130_fd_sc_hd__a2bb2o_4
X_23958_ _23949_/CLK _23958_/D HRESETn VGND VGND VPWR VPWR _17498_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22741__A1 _22539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13711_ _14072_/A VGND VGND VPWR VPWR _13711_/X sky130_fd_sc_hd__buf_2
XFILLER_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15759__B1 _24455_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22909_ _22968_/A _22909_/B VGND VGND VPWR VPWR _22909_/X sky130_fd_sc_hd__and2_4
X_14691_ _14682_/X _14690_/Y _14640_/X _14064_/Y _14643_/A VGND VGND VPWR VPWR _14692_/A
+ sky130_fd_sc_hd__a32o_4
X_23889_ _24962_/CLK _23889_/D HRESETn VGND VGND VPWR VPWR _18100_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22884__B _22884_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16430_ _24207_/Q VGND VGND VPWR VPWR _16430_/Y sky130_fd_sc_hd__inv_2
X_13642_ _13641_/Y _13639_/X _13398_/X _13639_/X VGND VGND VPWR VPWR _13642_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24813__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24886__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23061__A _20739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16361_ _24232_/Q VGND VGND VPWR VPWR _16361_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15779__A _15746_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _11667_/Y _13568_/X _13572_/X _13568_/B VGND VGND VPWR VPWR _13574_/A sky130_fd_sc_hd__o22a_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18100_ _18100_/A VGND VGND VPWR VPWR _21648_/A sky130_fd_sc_hd__inv_2
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15312_ _13613_/A _15310_/X HADDR[4] _15310_/X VGND VGND VPWR VPWR _24617_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ _12503_/X VGND VGND VPWR VPWR _12525_/B sky130_fd_sc_hd__inv_2
X_19080_ _19077_/Y _19079_/X _19059_/X _19079_/X VGND VGND VPWR VPWR _23462_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _14926_/Y _16286_/X _16291_/X _16286_/X VGND VGND VPWR VPWR _16292_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15526__A3 _15432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18031_ _19530_/A _18031_/B _18031_/C VGND VGND VPWR VPWR _19595_/A sky130_fd_sc_hd__or3_4
X_15243_ _15237_/X _15251_/B VGND VGND VPWR VPWR _15243_/X sky130_fd_sc_hd__or2_4
XANTENNA__13299__A _13299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12455_ _12454_/X VGND VGND VPWR VPWR _12455_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15174_ _15177_/A _15177_/B VGND VGND VPWR VPWR _15178_/B sky130_fd_sc_hd__or2_4
X_12386_ _25092_/Q _12384_/Y _12385_/Y _12382_/A VGND VGND VPWR VPWR _12387_/D sky130_fd_sc_hd__a2bb2o_4
X_14125_ _13492_/X VGND VGND VPWR VPWR _14126_/A sky130_fd_sc_hd__inv_2
XFILLER_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19982_ _19982_/A VGND VGND VPWR VPWR _19982_/X sky130_fd_sc_hd__buf_2
XFILLER_10_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12931__A _12922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14498__B1 _14484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14056_ _14055_/Y _14053_/X _13632_/X _14053_/X VGND VGND VPWR VPWR _14056_/X sky130_fd_sc_hd__a2bb2o_4
X_18933_ _18931_/Y _18927_/X _18932_/X _18927_/X VGND VGND VPWR VPWR _23514_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13007_ _25005_/Q _13007_/B VGND VGND VPWR VPWR _13008_/C sky130_fd_sc_hd__or2_4
XFILLER_136_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15019__A _15019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_29_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18864_ _18863_/Y _18859_/X _18795_/X _18859_/X VGND VGND VPWR VPWR _18864_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17815_ _17815_/A _17815_/B _17815_/C VGND VGND VPWR VPWR _17815_/X sky130_fd_sc_hd__or3_4
X_18795_ _18678_/X VGND VGND VPWR VPWR _18795_/X sky130_fd_sc_hd__buf_2
XANTENNA__15998__B1 _15801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17746_ _17894_/A _17746_/B _17746_/C VGND VGND VPWR VPWR _17746_/X sky130_fd_sc_hd__and3_4
X_14958_ _24275_/Q VGND VGND VPWR VPWR _14958_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21535__A2 _21533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13909_ _13845_/A _13908_/X _13905_/X _24904_/Q _13903_/X VGND VGND VPWR VPWR _13909_/X
+ sky130_fd_sc_hd__a32o_4
X_17677_ _17697_/A _17677_/B VGND VGND VPWR VPWR _17679_/B sky130_fd_sc_hd__or2_4
X_14889_ _14969_/A _14887_/Y _14888_/Y _14901_/A VGND VGND VPWR VPWR _14889_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16628_ _16628_/A VGND VGND VPWR VPWR _16632_/A sky130_fd_sc_hd__buf_2
X_19416_ _18068_/X _11761_/A _18666_/C VGND VGND VPWR VPWR _19417_/A sky130_fd_sc_hd__or3_4
XFILLER_56_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21299__A1 _21300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22375__A2_N _22372_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16559_ _16559_/A _16235_/B VGND VGND VPWR VPWR _16559_/X sky130_fd_sc_hd__or2_4
X_19347_ _13017_/B VGND VGND VPWR VPWR _19347_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22496__B1 _22482_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24556__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19278_ _21251_/A _19274_/X _19207_/X _19274_/X VGND VGND VPWR VPWR _19278_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16175__B1 _15777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18229_ _18223_/A _18223_/B _18225_/B _18228_/X VGND VGND VPWR VPWR _18229_/X sky130_fd_sc_hd__a211o_4
X_21240_ _21393_/A _19834_/Y VGND VGND VPWR VPWR _21240_/X sky130_fd_sc_hd__or2_4
XFILLER_116_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19664__B2 _19646_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21171_ _21130_/X _21171_/B _21171_/C VGND VGND VPWR VPWR _21171_/X sky130_fd_sc_hd__and3_4
XFILLER_102_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22034__B _21860_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20122_ _23082_/Q VGND VGND VPWR VPWR _20122_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20053_ _20983_/B _20048_/X _19755_/X _20035_/Y VGND VGND VPWR VPWR _20053_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19624__A _19636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24930_ _24928_/CLK _24930_/D HRESETn VGND VGND VPWR VPWR _13428_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_112_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23791__D MSI_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24861_ _23657_/CLK _14082_/X HRESETn VGND VGND VPWR VPWR _14081_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14768__A _24699_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23812_ _23824_/CLK _23812_/D HRESETn VGND VGND VPWR VPWR pwm_S7 sky130_fd_sc_hd__dfrtp_4
X_24792_ _24859_/CLK _24792_/D HRESETn VGND VGND VPWR VPWR _24792_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_39_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13464__B2 _13463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_192_0_HCLK clkbuf_7_96_0_HCLK/X VGND VGND VPWR VPWR _24405_/CLK sky130_fd_sc_hd__clkbuf_1
X_23743_ _23744_/CLK _23743_/D HRESETn VGND VGND VPWR VPWR _20635_/C sky130_fd_sc_hd__dfrtp_4
X_20955_ _20948_/X _20953_/X _22105_/A VGND VGND VPWR VPWR _20955_/X sky130_fd_sc_hd__o21a_4
XPHY_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_49_0_HCLK clkbuf_7_24_0_HCLK/X VGND VGND VPWR VPWR _25194_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_41_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23674_ _23680_/CLK _20380_/Y HRESETn VGND VGND VPWR VPWR _23674_/Q sky130_fd_sc_hd__dfrtp_4
X_20886_ _20886_/A _11725_/X VGND VGND VPWR VPWR _20886_/Y sky130_fd_sc_hd__nand2_4
XPHY_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22625_ _22011_/X _22623_/X _22322_/X _22624_/X VGND VGND VPWR VPWR _22625_/X sky130_fd_sc_hd__o22a_4
XPHY_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24297__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21113__B _21113_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16166__B1 _15855_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22556_ _16992_/A _22956_/B VGND VGND VPWR VPWR _22562_/B sky130_fd_sc_hd__or2_4
XANTENNA__15508__A3 _15507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12735__B _12638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24226__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21507_ _21376_/A _21505_/X _21506_/X VGND VGND VPWR VPWR _21507_/X sky130_fd_sc_hd__and3_4
XFILLER_33_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22487_ _22487_/A _22188_/X VGND VGND VPWR VPWR _22487_/X sky130_fd_sc_hd__and2_4
XANTENNA__19104__B1 _19038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12240_ _12094_/Y _12245_/B _12195_/X VGND VGND VPWR VPWR _12240_/Y sky130_fd_sc_hd__a21oi_4
X_24226_ _24225_/CLK _24226_/D HRESETn VGND VGND VPWR VPWR _16378_/A sky130_fd_sc_hd__dfrtp_4
X_21438_ _21570_/A _21438_/B _21437_/X VGND VGND VPWR VPWR _21457_/A sky130_fd_sc_hd__and3_4
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12171_ _12207_/A _12171_/B VGND VGND VPWR VPWR _12171_/X sky130_fd_sc_hd__or2_4
X_21369_ _21500_/A _21369_/B _21368_/X VGND VGND VPWR VPWR _21369_/X sky130_fd_sc_hd__and3_4
X_24157_ _24013_/CLK _24157_/D HRESETn VGND VGND VPWR VPWR _15099_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12751__A _12749_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16638__A1_N _14781_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23108_ _23085_/CLK _23108_/D VGND VGND VPWR VPWR _21649_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_1_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24088_ _24088_/CLK _24088_/D HRESETn VGND VGND VPWR VPWR _16774_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_89_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15930_ _15927_/Y _15923_/X _15753_/X _15929_/X VGND VGND VPWR VPWR _24389_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23861__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23039_ _23908_/Q _21651_/B _23037_/X _23038_/Y VGND VGND VPWR VPWR _23039_/X sky130_fd_sc_hd__a211o_4
XANTENNA__25085__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22962__A1 _22539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15861_ _15859_/Y _15854_/X _15772_/X _15860_/X VGND VGND VPWR VPWR _15861_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23056__A _20717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25014__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17600_ _16712_/Y _17603_/B _16748_/X VGND VGND VPWR VPWR _17600_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_67_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14812_ _14812_/A VGND VGND VPWR VPWR _14812_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18580_ _16354_/A _18517_/A _16354_/Y _18518_/A VGND VGND VPWR VPWR _18581_/D sky130_fd_sc_hd__o22a_4
X_15792_ _12800_/Y _15787_/X _15513_/X _15791_/X VGND VGND VPWR VPWR _24437_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22714__A1 _16692_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17531_ _17531_/A VGND VGND VPWR VPWR _23968_/D sky130_fd_sc_hd__inv_2
X_14743_ _14742_/Y VGND VGND VPWR VPWR _14743_/X sky130_fd_sc_hd__buf_2
X_11955_ _16301_/A _11954_/X VGND VGND VPWR VPWR _11955_/X sky130_fd_sc_hd__or2_4
XFILLER_45_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17462_ _17461_/X VGND VGND VPWR VPWR _17462_/Y sky130_fd_sc_hd__inv_2
X_14674_ _14640_/X _14673_/X _14055_/A _14643_/A VGND VGND VPWR VPWR _14674_/Y sky130_fd_sc_hd__a22oi_4
X_11886_ _11884_/A _11884_/B _11885_/Y VGND VGND VPWR VPWR _11886_/X sky130_fd_sc_hd__o21a_4
XFILLER_33_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15747__A3 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16413_ _16413_/A VGND VGND VPWR VPWR _16413_/Y sky130_fd_sc_hd__inv_2
X_19201_ _18678_/X VGND VGND VPWR VPWR _19201_/X sky130_fd_sc_hd__buf_2
X_13625_ _13624_/Y VGND VGND VPWR VPWR _13630_/C sky130_fd_sc_hd__buf_2
X_17393_ _17380_/X VGND VGND VPWR VPWR _17393_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12926__A _12925_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19132_ _17808_/B VGND VGND VPWR VPWR _19132_/Y sky130_fd_sc_hd__inv_2
X_16344_ _16343_/Y _16339_/X _16266_/X _16339_/X VGND VGND VPWR VPWR _16344_/X sky130_fd_sc_hd__a2bb2o_4
X_13556_ _11663_/Y _13555_/X VGND VGND VPWR VPWR _13557_/B sky130_fd_sc_hd__or2_4
XFILLER_73_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20101__A2_N _20098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12507_ _25081_/Q _12507_/B VGND VGND VPWR VPWR _12507_/X sky130_fd_sc_hd__or2_4
X_19063_ _17774_/B VGND VGND VPWR VPWR _19063_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16275_ _16268_/X _16269_/X _15505_/X _24267_/Q _16270_/X VGND VGND VPWR VPWR _16275_/X
+ sky130_fd_sc_hd__a32o_4
X_13487_ _13486_/Y _13482_/Y _13468_/A _13480_/X VGND VGND VPWR VPWR _24969_/D sky130_fd_sc_hd__o22a_4
XFILLER_51_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18014_ _18013_/Y _18008_/X _16617_/X _18007_/Y VGND VGND VPWR VPWR _18014_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15226_ _15226_/A _15225_/X _15226_/C VGND VGND VPWR VPWR _24653_/D sky130_fd_sc_hd__and3_4
X_12438_ _12438_/A VGND VGND VPWR VPWR _12444_/B sky130_fd_sc_hd__inv_2
XANTENNA__21453__A1 _17487_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15157_ _15156_/X VGND VGND VPWR VPWR _24672_/D sky130_fd_sc_hd__inv_2
XANTENNA__23949__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12369_ _25093_/Q VGND VGND VPWR VPWR _12415_/A sky130_fd_sc_hd__inv_2
XFILLER_113_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14108_ _14108_/A VGND VGND VPWR VPWR _14108_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21974__A _22629_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15088_ _14791_/X _15087_/X _14984_/X VGND VGND VPWR VPWR _15088_/Y sky130_fd_sc_hd__a21oi_4
X_19965_ _23143_/Q VGND VGND VPWR VPWR _19965_/Y sky130_fd_sc_hd__inv_2
X_14039_ _24874_/Q VGND VGND VPWR VPWR _14039_/Y sky130_fd_sc_hd__inv_2
X_18916_ _18915_/Y _18913_/X _18802_/X _18913_/X VGND VGND VPWR VPWR _23520_/D sky130_fd_sc_hd__a2bb2o_4
X_19896_ _23169_/Q VGND VGND VPWR VPWR _21382_/B sky130_fd_sc_hd__inv_2
XFILLER_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18082__B1 _13011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18847_ _23544_/Q VGND VGND VPWR VPWR _21211_/B sky130_fd_sc_hd__inv_2
XFILLER_95_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18778_ _17924_/B VGND VGND VPWR VPWR _18778_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18909__B1 _18817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_202_0_HCLK clkbuf_8_203_0_HCLK/A VGND VGND VPWR VPWR _24037_/CLK sky130_fd_sc_hd__clkbuf_1
X_17729_ _17729_/A VGND VGND VPWR VPWR _17817_/A sky130_fd_sc_hd__buf_2
XFILLER_36_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22181__A2 _22177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24737__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_8_0_HCLK clkbuf_7_4_0_HCLK/X VGND VGND VPWR VPWR _23292_/CLK sky130_fd_sc_hd__clkbuf_1
X_20740_ _20740_/A _20740_/B VGND VGND VPWR VPWR _20740_/X sky130_fd_sc_hd__and2_4
XFILLER_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21214__A _21214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20671_ _20671_/A VGND VGND VPWR VPWR _23754_/D sky130_fd_sc_hd__inv_2
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24390__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22410_ _22322_/X _22408_/X _22280_/X _22409_/X VGND VGND VPWR VPWR _22411_/B sky130_fd_sc_hd__o22a_4
XANTENNA__16148__B1 _15837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21141__B1 _18049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23390_ _23388_/CLK _23390_/D VGND VGND VPWR VPWR _23390_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22341_ _22691_/A _22341_/B _22341_/C VGND VGND VPWR VPWR _22381_/A sky130_fd_sc_hd__and3_4
XANTENNA__21692__A1 _16042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21692__B2 _22616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21868__B _21868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18523__A _18485_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22272_ _22272_/A _21357_/X VGND VGND VPWR VPWR _22272_/X sky130_fd_sc_hd__and2_4
X_25060_ _25050_/CLK _25060_/D HRESETn VGND VGND VPWR VPWR _12605_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22045__A _21490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21223_ _21383_/A _21223_/B VGND VGND VPWR VPWR _21223_/X sky130_fd_sc_hd__or2_4
XFILLER_105_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13382__B1 _13330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24011_ _24017_/CLK _17223_/X HRESETn VGND VGND VPWR VPWR _20735_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17139__A _17129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21444__B2 _21113_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16043__A _16043_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21154_ _21159_/A _21154_/B VGND VGND VPWR VPWR _21154_/X sky130_fd_sc_hd__or2_4
XANTENNA__23619__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24356__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20105_ _20105_/A VGND VGND VPWR VPWR _21621_/B sky130_fd_sc_hd__inv_2
XFILLER_67_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15882__A _24405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21085_ _14062_/Y _21083_/X _15288_/A _21425_/B VGND VGND VPWR VPWR _21090_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21747__A2 _21082_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20036_ _20035_/Y VGND VGND VPWR VPWR _20036_/X sky130_fd_sc_hd__buf_2
X_24913_ _23661_/CLK _13800_/X HRESETn VGND VGND VPWR VPWR scl_oen_o_S5 sky130_fd_sc_hd__dfstp_4
Xclkbuf_6_12_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_12_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16623__A1 _15619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16623__B2 _16622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24844_ _24962_/CLK _24844_/D HRESETn VGND VGND VPWR VPWR _24844_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24775_ _24776_/CLK _14341_/X HRESETn VGND VGND VPWR VPWR _21443_/A sky130_fd_sc_hd__dfrtp_4
X_21987_ _21292_/A VGND VGND VPWR VPWR _21987_/X sky130_fd_sc_hd__buf_2
XFILLER_57_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24478__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _23894_/Q VGND VGND VPWR VPWR _18065_/C sky130_fd_sc_hd__buf_2
XANTENNA__17602__A _16700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23726_ _24171_/CLK _23726_/D HRESETn VGND VGND VPWR VPWR _23726_/Q sky130_fd_sc_hd__dfrtp_4
X_20938_ _23025_/B _20935_/Y _22011_/A _20937_/X VGND VGND VPWR VPWR _20939_/B sky130_fd_sc_hd__a211o_4
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21380__B1 _21242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24407__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _23915_/Q VGND VGND VPWR VPWR _11671_/Y sky130_fd_sc_hd__inv_2
XPHY_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23657_ _23657_/CLK _20719_/X HRESETn VGND VGND VPWR VPWR _23657_/Q sky130_fd_sc_hd__dfrtp_4
X_20869_ _14009_/A _20844_/B VGND VGND VPWR VPWR _20869_/X sky130_fd_sc_hd__and2_4
XPHY_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _13408_/Y _14377_/A _22214_/A _24762_/Q VGND VGND VPWR VPWR _13418_/A sky130_fd_sc_hd__a2bb2o_4
XPHY_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16139__B1 _15828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22608_ _13334_/X VGND VGND VPWR VPWR _22608_/X sky130_fd_sc_hd__buf_2
X_14390_ _14387_/A _14386_/Y _14387_/C _14390_/D VGND VGND VPWR VPWR _14390_/X sky130_fd_sc_hd__and4_4
XPHY_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23588_ _23128_/CLK _23588_/D VGND VGND VPWR VPWR _17782_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_10_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24060__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13341_ _13341_/A VGND VGND VPWR VPWR _13341_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22539_ _21248_/X VGND VGND VPWR VPWR _22539_/X sky130_fd_sc_hd__buf_2
XFILLER_6_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16060_ _16058_/Y _16059_/X _11545_/X _16059_/X VGND VGND VPWR VPWR _16060_/X sky130_fd_sc_hd__a2bb2o_4
X_13272_ _13155_/X _13264_/X _13272_/C VGND VGND VPWR VPWR _13272_/X sky130_fd_sc_hd__and3_4
X_15011_ _15011_/A VGND VGND VPWR VPWR _15011_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13373__B1 _11626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12223_ _12190_/A _12219_/B _12222_/X VGND VGND VPWR VPWR _12223_/X sky130_fd_sc_hd__and3_4
X_24209_ _24262_/CLK _24209_/D HRESETn VGND VGND VPWR VPWR _24209_/Q sky130_fd_sc_hd__dfrtp_4
X_25189_ _23353_/CLK _25189_/D HRESETn VGND VGND VPWR VPWR _11701_/C sky130_fd_sc_hd__dfrtp_4
XANTENNA__21794__A _21292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12154_ _12154_/A VGND VGND VPWR VPWR _12154_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16311__B1 _16141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19750_ _19737_/Y VGND VGND VPWR VPWR _19750_/X sky130_fd_sc_hd__buf_2
X_12085_ _24555_/Q VGND VGND VPWR VPWR _12085_/Y sky130_fd_sc_hd__inv_2
X_16962_ _16202_/A _17034_/C _16149_/Y _24054_/Q VGND VGND VPWR VPWR _16962_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22935__A1 _21864_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18701_ _18699_/Y _18697_/X _18700_/X _18697_/X VGND VGND VPWR VPWR _18701_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15913_ _15916_/A _15418_/A VGND VGND VPWR VPWR _15913_/X sky130_fd_sc_hd__or2_4
X_16893_ _16825_/Y _16885_/B VGND VGND VPWR VPWR _16893_/X sky130_fd_sc_hd__or2_4
X_19681_ _19679_/Y _19680_/X _19614_/X _19680_/X VGND VGND VPWR VPWR _19681_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16614__A1 _15657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14840__A2_N _14838_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15844_ _24420_/Q VGND VGND VPWR VPWR _15844_/Y sky130_fd_sc_hd__inv_2
X_18632_ _20717_/A VGND VGND VPWR VPWR _18632_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15775_ HWDATA[18] VGND VGND VPWR VPWR _15775_/X sky130_fd_sc_hd__buf_2
X_18563_ _16349_/Y _18509_/A _16349_/Y _18509_/A VGND VGND VPWR VPWR _18566_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12987_ _12984_/A _12984_/B VGND VGND VPWR VPWR _12987_/Y sky130_fd_sc_hd__nand2_4
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24830__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14726_ _14726_/A VGND VGND VPWR VPWR _14726_/Y sky130_fd_sc_hd__inv_2
X_17514_ _17513_/X VGND VGND VPWR VPWR _17514_/Y sky130_fd_sc_hd__inv_2
X_11938_ _11938_/A _21300_/B VGND VGND VPWR VPWR _11939_/A sky130_fd_sc_hd__and2_4
X_18494_ _18494_/A VGND VGND VPWR VPWR _23833_/D sky130_fd_sc_hd__inv_2
XANTENNA__22775__D _22775_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24148__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17445_ _17445_/A VGND VGND VPWR VPWR _23978_/D sky130_fd_sc_hd__inv_2
XANTENNA__21034__A _21033_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14657_ _14643_/A VGND VGND VPWR VPWR _14657_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_32_0_HCLK clkbuf_8_33_0_HCLK/A VGND VGND VPWR VPWR _23112_/CLK sky130_fd_sc_hd__clkbuf_1
X_11869_ _11648_/X _11868_/Y _11866_/X VGND VGND VPWR VPWR _11869_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_33_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_95_0_HCLK clkbuf_8_95_0_HCLK/A VGND VGND VPWR VPWR _24723_/CLK sky130_fd_sc_hd__clkbuf_1
X_13608_ _14403_/A VGND VGND VPWR VPWR _13608_/X sky130_fd_sc_hd__buf_2
XANTENNA__12859__A1_N _12858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17376_ _17246_/Y _17373_/X VGND VGND VPWR VPWR _17376_/X sky130_fd_sc_hd__or2_4
XFILLER_20_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21969__A _21062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14588_ _14596_/A _14587_/X VGND VGND VPWR VPWR _14589_/B sky130_fd_sc_hd__or2_4
X_16327_ _16325_/Y _16321_/X _16251_/X _16326_/X VGND VGND VPWR VPWR _16327_/X sky130_fd_sc_hd__a2bb2o_4
X_19115_ _11635_/A VGND VGND VPWR VPWR _19115_/X sky130_fd_sc_hd__buf_2
X_13539_ _23752_/Q _23751_/Q _23753_/Q _20660_/B VGND VGND VPWR VPWR _13539_/X sky130_fd_sc_hd__or4_4
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22871__B1 _22530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19046_ _13212_/B VGND VGND VPWR VPWR _19046_/Y sky130_fd_sc_hd__inv_2
X_16258_ _14900_/Y _16257_/X _15855_/X _16257_/X VGND VGND VPWR VPWR _24276_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16550__B1 _16211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15209_ _15192_/A _15203_/B _15208_/Y VGND VGND VPWR VPWR _15209_/X sky130_fd_sc_hd__and3_4
XANTENNA__13364__B1 _11604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21426__A1 _22610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23783__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16189_ _16188_/Y _16184_/X _16096_/X _16184_/X VGND VGND VPWR VPWR _24301_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23712__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19948_ _19960_/A VGND VGND VPWR VPWR _19948_/X sky130_fd_sc_hd__buf_2
XANTENNA__22926__A1 _24153_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24989__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21209__A _21374_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19879_ _19878_/Y _19876_/X _19835_/X _19876_/X VGND VGND VPWR VPWR _23176_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14808__A2_N _24128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24918__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21910_ _21913_/A _21910_/B VGND VGND VPWR VPWR _21910_/X sky130_fd_sc_hd__or2_4
X_22890_ _22681_/A _22890_/B VGND VGND VPWR VPWR _22890_/X sky130_fd_sc_hd__and2_4
XFILLER_23_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21841_ _15456_/X VGND VGND VPWR VPWR _22178_/A sky130_fd_sc_hd__buf_2
XFILLER_71_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24571__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24560_ _24573_/CLK _24560_/D HRESETn VGND VGND VPWR VPWR _24560_/Q sky130_fd_sc_hd__dfrtp_4
X_21772_ _14443_/B VGND VGND VPWR VPWR _21777_/A sky130_fd_sc_hd__buf_2
XFILLER_63_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24500__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23511_ _23511_/CLK _18941_/X VGND VGND VPWR VPWR _17966_/B sky130_fd_sc_hd__dfxtp_4
X_20723_ _20723_/A _20723_/B VGND VGND VPWR VPWR _20723_/X sky130_fd_sc_hd__and2_4
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24491_ _25090_/CLK _15674_/X HRESETn VGND VGND VPWR VPWR _24491_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22982__B _22982_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23442_ _23442_/CLK _19135_/X VGND VGND VPWR VPWR _17846_/B sky130_fd_sc_hd__dfxtp_4
X_20654_ _23749_/Q _20649_/X _20653_/Y VGND VGND VPWR VPWR _20654_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20783__A _20751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_3_0_HCLK clkbuf_5_2_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__11602__B1 _25200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15877__A _24407_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20585_ _13533_/A _13533_/B VGND VGND VPWR VPWR _20585_/X sky130_fd_sc_hd__or2_4
X_23373_ _23374_/CLK _23373_/D VGND VGND VPWR VPWR _23373_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_104_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25112_ _25112_/CLK _25112_/D HRESETn VGND VGND VPWR VPWR _12177_/A sky130_fd_sc_hd__dfrtp_4
X_22324_ _16527_/Y _22488_/B VGND VGND VPWR VPWR _22324_/X sky130_fd_sc_hd__and2_4
XFILLER_136_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13397__A _16302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25043_ _25046_/CLK _12756_/X HRESETn VGND VGND VPWR VPWR _25043_/Q sky130_fd_sc_hd__dfrtp_4
X_22255_ _22852_/A VGND VGND VPWR VPWR _22256_/B sky130_fd_sc_hd__buf_2
XFILLER_117_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21968__A2 _21923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21206_ _21371_/A _19941_/Y VGND VGND VPWR VPWR _21207_/C sky130_fd_sc_hd__or2_4
X_22186_ _21569_/A _22185_/X VGND VGND VPWR VPWR _22201_/B sky130_fd_sc_hd__and2_4
X_21137_ _21469_/A _19548_/Y VGND VGND VPWR VPWR _21140_/B sky130_fd_sc_hd__or2_4
XFILLER_28_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22917__A1 _16621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22917__B2 _21694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18046__B1 _21335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21068_ _20926_/A VGND VGND VPWR VPWR _22322_/A sky130_fd_sc_hd__buf_2
XFILLER_115_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21119__A _11952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12330__A1 _12328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24659__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12910_ _12921_/A _12910_/B _12910_/C VGND VGND VPWR VPWR _12910_/X sky130_fd_sc_hd__and3_4
X_20019_ _20019_/A VGND VGND VPWR VPWR _21809_/B sky130_fd_sc_hd__inv_2
XFILLER_24_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12330__B2 _12329_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13890_ _13890_/A VGND VGND VPWR VPWR _13891_/A sky130_fd_sc_hd__buf_2
XFILLER_46_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14021__A _16301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12841_ _12947_/A _24446_/Q _22712_/A _12790_/Y VGND VGND VPWR VPWR _12844_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24827_ _24824_/CLK _24827_/D HRESETn VGND VGND VPWR VPWR _24827_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_76_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17245__A1_N _25200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15280__B1 _15279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15560_ _15557_/Y _15558_/X _15559_/X _15558_/X VGND VGND VPWR VPWR _15560_/X sky130_fd_sc_hd__a2bb2o_4
X_12772_ _12651_/D _12663_/B _12674_/X _12770_/B VGND VGND VPWR VPWR _12773_/A sky130_fd_sc_hd__a211o_4
XPHY_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24758_ _24928_/CLK _24758_/D HRESETn VGND VGND VPWR VPWR _14414_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24241__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14511_/A VGND VGND VPWR VPWR _21756_/A sky130_fd_sc_hd__inv_2
XFILLER_76_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _13612_/A _12060_/A VGND VGND VPWR VPWR _11723_/X sky130_fd_sc_hd__and2_4
XPHY_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23709_ _24612_/CLK _20483_/X HRESETn VGND VGND VPWR VPWR _13509_/B sky130_fd_sc_hd__dfrtp_4
X_15491_ _12095_/Y _15487_/X _11566_/X _15490_/X VGND VGND VPWR VPWR _15491_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11841__B1 _11839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_19_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24689_ _24264_/CLK _24689_/D HRESETn VGND VGND VPWR VPWR _24689_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _23896_/Q _17227_/B _17228_/Y VGND VGND VPWR VPWR _17230_/X sky130_fd_sc_hd__o21a_4
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _21012_/A VGND VGND VPWR VPWR _14443_/B sky130_fd_sc_hd__buf_2
XFILLER_120_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _13571_/A _23922_/Q _13571_/A _23922_/Q VGND VGND VPWR VPWR _11654_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17161_ _17161_/A _17161_/B VGND VGND VPWR VPWR _17161_/X sky130_fd_sc_hd__or2_4
XANTENNA__15787__A _15767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14373_ _14424_/A _13442_/A VGND VGND VPWR VPWR _14373_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__19259__A _16043_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11585_ _11585_/A VGND VGND VPWR VPWR _11585_/X sky130_fd_sc_hd__buf_2
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16112_ _16084_/A VGND VGND VPWR VPWR _16112_/X sky130_fd_sc_hd__buf_2
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13324_ _11950_/X _14195_/B _22510_/B VGND VGND VPWR VPWR _13324_/X sky130_fd_sc_hd__or3_4
XFILLER_70_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17092_ _17074_/A _17092_/B _17092_/C VGND VGND VPWR VPWR _17093_/A sky130_fd_sc_hd__or3_4
XFILLER_13_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17875__A3 _17874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16043_ _16043_/A _23763_/Q _16041_/X _22265_/B VGND VGND VPWR VPWR _16043_/X sky130_fd_sc_hd__and4_4
X_13255_ _11735_/Y _13247_/X _13254_/X VGND VGND VPWR VPWR _13255_/X sky130_fd_sc_hd__and3_4
XFILLER_100_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12206_ _12167_/Y _12183_/B _12171_/B _12183_/A VGND VGND VPWR VPWR _12207_/B sky130_fd_sc_hd__or4_4
XFILLER_135_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13186_ _11741_/X VGND VGND VPWR VPWR _13219_/A sky130_fd_sc_hd__buf_2
X_19802_ _19802_/A VGND VGND VPWR VPWR _19802_/X sky130_fd_sc_hd__buf_2
X_12137_ _12174_/B _24562_/Q _12172_/A _12088_/Y VGND VGND VPWR VPWR _12137_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17507__A _23012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17994_ _17982_/X _17990_/X _17993_/X _23917_/Q _17983_/X VGND VGND VPWR VPWR _17994_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_46_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22908__A1 _15463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22908__B2 _22576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19733_ _19733_/A VGND VGND VPWR VPWR _19733_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21029__A _20814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12068_ SSn_S3 _12067_/Y _11981_/X _12067_/Y VGND VGND VPWR VPWR _25135_/D sky130_fd_sc_hd__a2bb2o_4
X_16945_ _16922_/A _16922_/B _16942_/Y _16858_/X VGND VGND VPWR VPWR _16946_/A sky130_fd_sc_hd__a211o_4
XFILLER_49_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11555__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19664_ _20984_/B _19659_/X _19641_/X _19646_/Y VGND VGND VPWR VPWR _23255_/D sky130_fd_sc_hd__a2bb2o_4
X_16876_ _16876_/A VGND VGND VPWR VPWR _16881_/B sky130_fd_sc_hd__inv_2
XANTENNA__16599__B1 _15501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24329__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18615_ _18615_/A _18614_/X VGND VGND VPWR VPWR _18616_/B sky130_fd_sc_hd__or2_4
X_15827_ _15826_/X VGND VGND VPWR VPWR _15827_/X sky130_fd_sc_hd__buf_2
XFILLER_20_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19595_ _19595_/A VGND VGND VPWR VPWR _19613_/A sky130_fd_sc_hd__inv_2
XANTENNA__19537__B1 _11839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15758_ _12791_/Y _15752_/X _15756_/X _15757_/X VGND VGND VPWR VPWR _15758_/X sky130_fd_sc_hd__a2bb2o_4
X_18546_ _23818_/Q _18546_/B VGND VGND VPWR VPWR _18547_/C sky130_fd_sc_hd__or2_4
XFILLER_33_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14709_ _14709_/A VGND VGND VPWR VPWR _14709_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11832__B1 RsRx_S1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15689_ _15689_/A VGND VGND VPWR VPWR _15689_/X sky130_fd_sc_hd__buf_2
X_18477_ _18476_/X VGND VGND VPWR VPWR _23837_/D sky130_fd_sc_hd__inv_2
XFILLER_61_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17428_ _17412_/B _17426_/Y _17428_/C VGND VGND VPWR VPWR _23984_/D sky130_fd_sc_hd__and3_4
XFILLER_127_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23964__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17359_ _17306_/Y _17362_/B _17336_/X VGND VGND VPWR VPWR _17359_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__25188__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20370_ _14045_/Y _20367_/X _20358_/X _20369_/X VGND VGND VPWR VPWR _20371_/A sky130_fd_sc_hd__a211o_4
XANTENNA__25117__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19029_ _19029_/A VGND VGND VPWR VPWR _20998_/B sky130_fd_sc_hd__inv_2
XANTENNA__18801__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22040_ _22146_/B _22029_/X _22033_/Y _21080_/Y _22039_/X VGND VGND VPWR VPWR _22040_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_133_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16321__A _16339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23991_ _24005_/CLK _17404_/X HRESETn VGND VGND VPWR VPWR _17315_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_60_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22942_ _21540_/X _22940_/X _20839_/X _22941_/X VGND VGND VPWR VPWR _22942_/X sky130_fd_sc_hd__o22a_4
XFILLER_112_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20778__A _20778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22873_ _22872_/X VGND VGND VPWR VPWR _22873_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24612_ _24612_/CLK _15334_/X HRESETn VGND VGND VPWR VPWR _15331_/A sky130_fd_sc_hd__dfrtp_4
X_21824_ _21913_/A _21824_/B VGND VGND VPWR VPWR _21824_/X sky130_fd_sc_hd__or2_4
XFILLER_36_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17003__B2 _24042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24543_ _24618_/CLK _15530_/X HRESETn VGND VGND VPWR VPWR _20413_/A sky130_fd_sc_hd__dfrtp_4
X_21755_ _14500_/Y _23393_/Q _21756_/A _21756_/B VGND VGND VPWR VPWR _21755_/X sky130_fd_sc_hd__o22a_4
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20706_ _23808_/Q _20705_/B _23807_/Q _20705_/X VGND VGND VPWR VPWR _20706_/X sky130_fd_sc_hd__o22a_4
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24474_ _24307_/CLK _15700_/X HRESETn VGND VGND VPWR VPWR _24474_/Q sky130_fd_sc_hd__dfrtp_4
X_21686_ _21675_/A _21683_/X _21685_/X VGND VGND VPWR VPWR _21686_/X sky130_fd_sc_hd__and3_4
XANTENNA__16762__B1 _24422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23425_ _23425_/CLK _23425_/D VGND VGND VPWR VPWR _19181_/A sky130_fd_sc_hd__dfxtp_4
X_20637_ _20621_/X _20636_/X _24176_/Q _20624_/X VGND VGND VPWR VPWR _23745_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23634__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16514__B1 _16266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23356_ _23356_/CLK _23356_/D VGND VGND VPWR VPWR _13144_/B sky130_fd_sc_hd__dfxtp_4
X_20568_ _16548_/Y _20553_/X _20562_/X _20567_/X VGND VGND VPWR VPWR _20568_/X sky130_fd_sc_hd__o22a_4
X_22307_ _22307_/A _22256_/B VGND VGND VPWR VPWR _22307_/X sky130_fd_sc_hd__and2_4
XANTENNA__14016__A _14016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23287_ _23383_/CLK _19572_/X VGND VGND VPWR VPWR _23287_/Q sky130_fd_sc_hd__dfxtp_4
X_20499_ _20499_/A _20499_/B _20499_/C _20517_/A VGND VGND VPWR VPWR _20499_/X sky130_fd_sc_hd__or4_4
XANTENNA__18711__A _13644_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13040_ _11753_/A _13038_/X _13040_/C VGND VGND VPWR VPWR _13040_/X sky130_fd_sc_hd__and3_4
X_25026_ _24566_/CLK _12940_/X HRESETn VGND VGND VPWR VPWR _22712_/A sky130_fd_sc_hd__dfrtp_4
X_22238_ _20786_/A VGND VGND VPWR VPWR _22238_/X sky130_fd_sc_hd__buf_2
XANTENNA__12000__B1 _11620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12551__B2 _24527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22169_ _22952_/B VGND VGND VPWR VPWR _22175_/A sky130_fd_sc_hd__buf_2
XFILLER_117_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14828__B1 _15019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16231__A _16231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14991_ _15014_/A _14989_/X _14991_/C VGND VGND VPWR VPWR _14991_/X sky130_fd_sc_hd__and3_4
XFILLER_43_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24493__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13942_ _24887_/Q _13941_/X _24888_/Q VGND VGND VPWR VPWR _13943_/B sky130_fd_sc_hd__or3_4
X_16730_ _15963_/Y _22473_/A _15963_/Y _22473_/A VGND VGND VPWR VPWR _16730_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21574__B1 _21292_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24422__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16661_ _14709_/Y _16659_/X _15788_/A _16659_/X VGND VGND VPWR VPWR _16661_/X sky130_fd_sc_hd__a2bb2o_4
X_13873_ _13873_/A VGND VGND VPWR VPWR _13877_/C sky130_fd_sc_hd__inv_2
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15612_ _15585_/A VGND VGND VPWR VPWR _15612_/X sky130_fd_sc_hd__buf_2
X_18400_ _24212_/Q _18468_/A _16423_/Y _23833_/Q VGND VGND VPWR VPWR _18401_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12824_ _25010_/Q VGND VGND VPWR VPWR _21840_/A sky130_fd_sc_hd__inv_2
X_16592_ _14838_/Y _16587_/X _16266_/X _16587_/X VGND VGND VPWR VPWR _16592_/X sky130_fd_sc_hd__a2bb2o_4
X_19380_ _19380_/A VGND VGND VPWR VPWR _19380_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14810__A1_N _15003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15543_ _19821_/A VGND VGND VPWR VPWR _19448_/A sky130_fd_sc_hd__buf_2
X_18331_ _18327_/A _18327_/B VGND VGND VPWR VPWR _18332_/B sky130_fd_sc_hd__nand2_4
X_12755_ _12636_/X VGND VGND VPWR VPWR _12755_/X sky130_fd_sc_hd__buf_2
XFILLER_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _11706_/A VGND VGND VPWR VPWR _11707_/A sky130_fd_sc_hd__inv_2
X_18262_ _18262_/A VGND VGND VPWR VPWR _18284_/A sky130_fd_sc_hd__buf_2
XPHY_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _12144_/Y _15472_/X _15332_/X _15472_/X VGND VGND VPWR VPWR _15474_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12686_/A VGND VGND VPWR VPWR _12686_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ _14373_/Y _14424_/X _14371_/X _14415_/X _14424_/A VGND VGND VPWR VPWR _24754_/D
+ sky130_fd_sc_hd__a32o_4
X_17213_ _17213_/A VGND VGND VPWR VPWR _17213_/X sky130_fd_sc_hd__buf_2
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11637_ _11633_/Y _11521_/A _11636_/X _11521_/A VGND VGND VPWR VPWR _25192_/D sky130_fd_sc_hd__a2bb2o_4
X_18193_ _18485_/C VGND VGND VPWR VPWR _18468_/C sky130_fd_sc_hd__buf_2
XFILLER_50_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16406__A _24217_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_106_0_HCLK clkbuf_7_53_0_HCLK/X VGND VGND VPWR VPWR _24425_/CLK sky130_fd_sc_hd__clkbuf_1
X_17144_ _17144_/A _17153_/B VGND VGND VPWR VPWR _17145_/B sky130_fd_sc_hd__or2_4
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14356_ _14349_/Y _13900_/B _20179_/C VGND VGND VPWR VPWR _14356_/X sky130_fd_sc_hd__o21a_4
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11568_ _11568_/A VGND VGND VPWR VPWR _11568_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25210__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_169_0_HCLK clkbuf_7_84_0_HCLK/X VGND VGND VPWR VPWR _23313_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22841__A3 _22839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13307_ _13171_/A _13307_/B _13306_/X VGND VGND VPWR VPWR _13311_/B sky130_fd_sc_hd__and3_4
X_17075_ _17074_/X VGND VGND VPWR VPWR _17075_/Y sky130_fd_sc_hd__inv_2
X_14287_ _16559_/A _18633_/A VGND VGND VPWR VPWR _14288_/A sky130_fd_sc_hd__nor2_4
X_11499_ _11499_/A _12060_/A VGND VGND VPWR VPWR _14013_/B sky130_fd_sc_hd__or2_4
XFILLER_48_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16026_ _14573_/A _18759_/B _14573_/A _18759_/B VGND VGND VPWR VPWR _16680_/A sky130_fd_sc_hd__a2bb2o_4
X_13238_ _13238_/A _13238_/B _13237_/X VGND VGND VPWR VPWR _13239_/C sky130_fd_sc_hd__and3_4
XFILLER_48_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13169_ _13169_/A VGND VGND VPWR VPWR _13301_/A sky130_fd_sc_hd__buf_2
XFILLER_123_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16141__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14819__B1 _15087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23003__B1 _25221_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17977_ _17987_/A VGND VGND VPWR VPWR _17977_/X sky130_fd_sc_hd__buf_2
XFILLER_46_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15492__B1 _11570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19716_ _19716_/A VGND VGND VPWR VPWR _21808_/B sky130_fd_sc_hd__inv_2
XANTENNA__19452__A _19452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16928_ _16834_/D _16927_/X VGND VGND VPWR VPWR _16932_/B sky130_fd_sc_hd__or2_4
XFILLER_78_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20598__A _20647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24163__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19647_ _19646_/Y VGND VGND VPWR VPWR _19647_/X sky130_fd_sc_hd__buf_2
XFILLER_93_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16859_ _16853_/A _16853_/B _16858_/X _16854_/Y VGND VGND VPWR VPWR _16859_/X sky130_fd_sc_hd__a211o_4
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19578_ _23285_/Q VGND VGND VPWR VPWR _19578_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18529_ _18420_/Y _18529_/B VGND VGND VPWR VPWR _18530_/C sky130_fd_sc_hd__or2_4
XANTENNA__19930__B1 _19445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21540_ _22637_/A VGND VGND VPWR VPWR _21540_/X sky130_fd_sc_hd__buf_2
XANTENNA__20540__B2 _20465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21471_ _21147_/A _21471_/B _21470_/X VGND VGND VPWR VPWR _21471_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_65_0_HCLK clkbuf_6_32_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_65_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23210_ _23282_/CLK _23210_/D VGND VGND VPWR VPWR _23210_/Q sky130_fd_sc_hd__dfxtp_4
X_20422_ _13499_/A _21020_/A _13499_/Y VGND VGND VPWR VPWR _20422_/Y sky130_fd_sc_hd__a21oi_4
X_24190_ _24222_/CLK _24190_/D HRESETn VGND VGND VPWR VPWR _24190_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23141_ _23332_/CLK _23141_/D VGND VGND VPWR VPWR _23141_/Q sky130_fd_sc_hd__dfxtp_4
X_20353_ _17173_/A _17173_/B VGND VGND VPWR VPWR _20353_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__21876__B _15639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20284_ _14239_/Y _20273_/X _14266_/X _20283_/X VGND VGND VPWR VPWR _20285_/A sky130_fd_sc_hd__a211o_4
X_23072_ _23993_/CLK _23072_/D VGND VGND VPWR VPWR _23072_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_136_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12533__A1 _12389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24933__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22023_ _22223_/A _22007_/X _22010_/Y _22022_/Y VGND VGND VPWR VPWR _22023_/X sky130_fd_sc_hd__a211o_4
XANTENNA__19997__B1 _19424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_5_25_0_HCLK_A clkbuf_4_12_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15890__A _16369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23974_ _23898_/CLK _17475_/X HRESETn VGND VGND VPWR VPWR _21801_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__11639__A3 _13398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21556__B1 _14055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22925_ _14956_/A _22859_/X _22338_/A VGND VGND VPWR VPWR _22925_/X sky130_fd_sc_hd__o21a_4
XFILLER_44_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22856_ _22982_/A _22853_/X _22854_/X _22856_/D VGND VGND VPWR VPWR _22856_/X sky130_fd_sc_hd__or4_4
XANTENNA__15786__B2 _15746_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21807_ _20833_/X _21807_/B VGND VGND VPWR VPWR _21807_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__23886__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21859__B2 _20757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22787_ _20820_/X _22786_/X VGND VGND VPWR VPWR _22787_/Y sky130_fd_sc_hd__nor2_4
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18706__A _16291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19921__B1 _19835_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12540_ _20739_/A VGND VGND VPWR VPWR _12540_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23815__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24526_ _24523_/CLK _24526_/D HRESETn VGND VGND VPWR VPWR _24526_/Q sky130_fd_sc_hd__dfrtp_4
X_21738_ _21738_/A VGND VGND VPWR VPWR _21738_/Y sky130_fd_sc_hd__inv_2
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25039__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22228__A _22228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12471_ _12460_/A _12471_/B _12470_/X VGND VGND VPWR VPWR _25091_/D sky130_fd_sc_hd__and3_4
XANTENNA__22808__B1 _20780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24457_ _24502_/CLK _15755_/X HRESETn VGND VGND VPWR VPWR _22913_/A sky130_fd_sc_hd__dfrtp_4
X_21669_ _21677_/A _21669_/B VGND VGND VPWR VPWR _21669_/X sky130_fd_sc_hd__or2_4
X_14210_ _20235_/D _14200_/X _14209_/X _14202_/X VGND VGND VPWR VPWR _14210_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23408_ _23979_/CLK _19230_/X VGND VGND VPWR VPWR _23408_/Q sky130_fd_sc_hd__dfxtp_4
X_15190_ _15190_/A _15190_/B VGND VGND VPWR VPWR _15192_/B sky130_fd_sc_hd__or2_4
X_24388_ _24425_/CLK _15932_/X HRESETn VGND VGND VPWR VPWR _22910_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_137_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14141_ _24842_/Q _14120_/B _24841_/Q _14115_/X VGND VGND VPWR VPWR _14141_/X sky130_fd_sc_hd__o22a_4
XFILLER_126_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23339_ _23336_/CLK _23339_/D VGND VGND VPWR VPWR _13187_/B sky130_fd_sc_hd__dfxtp_4
X_14072_ _14072_/A _13791_/A VGND VGND VPWR VPWR _15236_/A sky130_fd_sc_hd__or2_4
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23059__A _20737_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13023_ _13042_/A _13023_/B VGND VGND VPWR VPWR _13024_/C sky130_fd_sc_hd__or2_4
X_17900_ _17796_/X _23521_/Q VGND VGND VPWR VPWR _17901_/C sky130_fd_sc_hd__or2_4
XANTENNA__24674__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25009_ _25009_/CLK _12997_/Y HRESETn VGND VGND VPWR VPWR _25009_/Q sky130_fd_sc_hd__dfrtp_4
X_18880_ _18739_/X VGND VGND VPWR VPWR _18880_/X sky130_fd_sc_hd__buf_2
XFILLER_121_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24603__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17831_ _17898_/A _17831_/B _17830_/X VGND VGND VPWR VPWR _17842_/B sky130_fd_sc_hd__or3_4
XFILLER_126_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15474__B1 _15332_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22339__A2 _22477_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17762_ _14569_/A _17759_/X _17761_/X VGND VGND VPWR VPWR _17762_/X sky130_fd_sc_hd__and3_4
X_14974_ _14974_/A _14973_/X VGND VGND VPWR VPWR _14974_/X sky130_fd_sc_hd__or2_4
XFILLER_94_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23000__A3 _22251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19501_ _19488_/Y VGND VGND VPWR VPWR _19501_/X sky130_fd_sc_hd__buf_2
X_16713_ _22192_/A _22202_/A _15977_/Y _16712_/Y VGND VGND VPWR VPWR _16716_/C sky130_fd_sc_hd__o22a_4
XFILLER_75_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13925_ _13925_/A _13925_/B _13925_/C _13925_/D VGND VGND VPWR VPWR _13926_/B sky130_fd_sc_hd__or4_4
X_17693_ _17697_/A _23470_/Q VGND VGND VPWR VPWR _17693_/X sky130_fd_sc_hd__or2_4
XFILLER_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19432_ _19417_/Y VGND VGND VPWR VPWR _19432_/X sky130_fd_sc_hd__buf_2
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13856_ _13824_/X _13825_/X _24905_/Q _24904_/Q VGND VGND VPWR VPWR _13856_/X sky130_fd_sc_hd__a211o_4
X_16644_ _14737_/Y _16639_/X _16261_/X _16643_/X VGND VGND VPWR VPWR _24112_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12807_ _22133_/A _22126_/A _12805_/Y _12806_/Y VGND VGND VPWR VPWR _12807_/X sky130_fd_sc_hd__o22a_4
X_19363_ _19349_/Y VGND VGND VPWR VPWR _19363_/X sky130_fd_sc_hd__buf_2
X_13787_ _13787_/A VGND VGND VPWR VPWR _13787_/Y sky130_fd_sc_hd__inv_2
X_16575_ _16575_/A VGND VGND VPWR VPWR _16584_/A sky130_fd_sc_hd__buf_2
XFILLER_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18314_ _18210_/B _18304_/X VGND VGND VPWR VPWR _18314_/Y sky130_fd_sc_hd__nand2_4
X_12738_ _12593_/Y _12737_/X VGND VGND VPWR VPWR _12739_/B sky130_fd_sc_hd__or2_4
X_15526_ _15503_/X _15504_/X _15432_/X _24545_/Q _15466_/A VGND VGND VPWR VPWR _15526_/X
+ sky130_fd_sc_hd__a32o_4
X_19294_ _19293_/Y _19289_/X _11853_/X _19289_/X VGND VGND VPWR VPWR _23386_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14764__A1_N _15019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22138__A _22023_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15457_ _15414_/A _15456_/X VGND VGND VPWR VPWR _15659_/B sky130_fd_sc_hd__or2_4
X_18245_ _18221_/A _18243_/A VGND VGND VPWR VPWR _18246_/C sky130_fd_sc_hd__or2_4
X_12669_ _12669_/A _12727_/A _12663_/A VGND VGND VPWR VPWR _12672_/B sky130_fd_sc_hd__or3_4
XFILLER_30_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14408_ _14383_/B _14399_/X _14407_/Y _14403_/X _13438_/A VGND VGND VPWR VPWR _14408_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21977__A _21050_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15388_ _22008_/A _15381_/X _15386_/X _15387_/X VGND VGND VPWR VPWR _24591_/D sky130_fd_sc_hd__a2bb2o_4
X_18176_ _22479_/A _23860_/Q _22479_/A _23860_/Q VGND VGND VPWR VPWR _18177_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20881__A _20881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14339_ _14335_/X _14338_/X _24788_/Q _14331_/X VGND VGND VPWR VPWR _14339_/X sky130_fd_sc_hd__o22a_4
X_17127_ _24040_/Q _17127_/B VGND VGND VPWR VPWR _17129_/B sky130_fd_sc_hd__or2_4
XFILLER_102_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21696__B _21251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17058_ _17021_/Y _17055_/X _17051_/B _17057_/X VGND VGND VPWR VPWR _17058_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22027__B2 _22218_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16009_ _15438_/A _15437_/X VGND VGND VPWR VPWR _16009_/X sky130_fd_sc_hd__or2_4
Xclkbuf_4_7_0_HCLK clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24344__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22601__A _21434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15480__A3 _15479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20971_ _20971_/A VGND VGND VPWR VPWR _20972_/A sky130_fd_sc_hd__buf_2
XFILLER_53_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15215__A _15158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22710_ _21030_/X _22709_/X _22646_/X _24416_/Q _22647_/X VGND VGND VPWR VPWR _22710_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_96_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23690_ _24728_/CLK _23690_/D HRESETn VGND VGND VPWR VPWR _23690_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16728__A2_N _17481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22641_ _21292_/A VGND VGND VPWR VPWR _22641_/X sky130_fd_sc_hd__buf_2
XFILLER_34_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22572_ _22572_/A _22567_/X _22572_/C VGND VGND VPWR VPWR _22572_/X sky130_fd_sc_hd__or3_4
XFILLER_90_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25132__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24311_ _24049_/CLK _24311_/D HRESETn VGND VGND VPWR VPWR _16162_/A sky130_fd_sc_hd__dfrtp_4
X_21523_ _21387_/A _21521_/X _21522_/X VGND VGND VPWR VPWR _21523_/X sky130_fd_sc_hd__and3_4
XFILLER_55_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24242_ _24262_/CLK _16337_/X HRESETn VGND VGND VPWR VPWR _24242_/Q sky130_fd_sc_hd__dfrtp_4
X_21454_ _12389_/X _15456_/X _21453_/X VGND VGND VPWR VPWR _21454_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22266__B2 _16305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16285__A1_N _14887_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20405_ _20405_/A _20212_/B VGND VGND VPWR VPWR _20405_/X sky130_fd_sc_hd__or2_4
XFILLER_119_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20816__A2 _22429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24173_ _24171_/CLK _16519_/X HRESETn VGND VGND VPWR VPWR _24173_/Q sky130_fd_sc_hd__dfrtp_4
X_21385_ _21385_/A _19522_/Y VGND VGND VPWR VPWR _21387_/B sky130_fd_sc_hd__or2_4
Xclkbuf_8_152_0_HCLK clkbuf_7_76_0_HCLK/X VGND VGND VPWR VPWR _25044_/CLK sky130_fd_sc_hd__clkbuf_1
X_23124_ _23100_/CLK _20018_/X VGND VGND VPWR VPWR _23124_/Q sky130_fd_sc_hd__dfxtp_4
X_20336_ _20336_/A _20179_/B VGND VGND VPWR VPWR _20336_/X sky130_fd_sc_hd__or2_4
XFILLER_66_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22569__A2 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23055_ _23042_/X VGND VGND VPWR VPWR IRQ[3] sky130_fd_sc_hd__buf_2
X_20267_ _20162_/X _20234_/X _20249_/B _14309_/X _20171_/B VGND VGND VPWR VPWR _23776_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_62_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24085__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22006_ _22006_/A _22006_/B VGND VGND VPWR VPWR _22006_/Y sky130_fd_sc_hd__nor2_4
X_20198_ _14204_/Y _14309_/X _20163_/C VGND VGND VPWR VPWR _20198_/X sky130_fd_sc_hd__a21o_4
XFILLER_27_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22511__A _22510_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24014__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11971_ _11965_/Y VGND VGND VPWR VPWR _11971_/X sky130_fd_sc_hd__buf_2
XFILLER_56_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23957_ _23957_/CLK _23957_/D HRESETn VGND VGND VPWR VPWR _22473_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12749__A _12749_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13710_ _23659_/Q VGND VGND VPWR VPWR _14072_/A sky130_fd_sc_hd__buf_2
XFILLER_5_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22908_ _15463_/X _22907_/X _22835_/X _24423_/Q _22576_/A VGND VGND VPWR VPWR _22909_/B
+ sky130_fd_sc_hd__a32o_4
X_14690_ _14681_/A _14633_/X VGND VGND VPWR VPWR _14690_/Y sky130_fd_sc_hd__nand2_4
X_23888_ _25186_/CLK _23888_/D HRESETn VGND VGND VPWR VPWR _18089_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20966__A _20966_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13641_ _24942_/Q VGND VGND VPWR VPWR _13641_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22839_ _22835_/A VGND VGND VPWR VPWR _22839_/X sky130_fd_sc_hd__buf_2
XFILLER_77_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16360_ _16358_/Y _16359_/X _16100_/X _16359_/X VGND VGND VPWR VPWR _16360_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ _13572_/A _13571_/X VGND VGND VPWR VPWR _13572_/X sky130_fd_sc_hd__or2_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15311_ _21581_/A _15310_/X HADDR[5] _15310_/X VGND VGND VPWR VPWR _15311_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _12509_/A _12511_/D _12523_/C VGND VGND VPWR VPWR _12523_/X sky130_fd_sc_hd__and3_4
XFILLER_38_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24509_ _25034_/CLK _24509_/D HRESETn VGND VGND VPWR VPWR _24509_/Q sky130_fd_sc_hd__dfrtp_4
X_16291_ _16291_/A VGND VGND VPWR VPWR _16291_/X sky130_fd_sc_hd__buf_2
XFILLER_13_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15242_ _15262_/A VGND VGND VPWR VPWR _15251_/B sky130_fd_sc_hd__buf_2
X_18030_ _18030_/A _17625_/A _18038_/A VGND VGND VPWR VPWR _18031_/C sky130_fd_sc_hd__or3_4
X_12454_ _12448_/A _12448_/B _12453_/X _12449_/Y VGND VGND VPWR VPWR _12454_/X sky130_fd_sc_hd__a211o_4
XFILLER_138_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24855__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15173_ _15179_/A _15183_/B VGND VGND VPWR VPWR _15177_/B sky130_fd_sc_hd__or2_4
XANTENNA__15795__A _15767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12385_ _22678_/A VGND VGND VPWR VPWR _12385_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14124_ _14124_/A VGND VGND VPWR VPWR _14124_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19981_ _19981_/A VGND VGND VPWR VPWR _21389_/B sky130_fd_sc_hd__inv_2
XANTENNA__18881__B1 _18880_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14498__B2 _14497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14055_ _14055_/A VGND VGND VPWR VPWR _14055_/Y sky130_fd_sc_hd__inv_2
X_18932_ _18678_/X VGND VGND VPWR VPWR _18932_/X sky130_fd_sc_hd__buf_2
XFILLER_10_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16806__A1_N _15830_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14204__A _24822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13006_ _12925_/X _12999_/X _13005_/Y VGND VGND VPWR VPWR _25006_/D sky130_fd_sc_hd__and3_4
X_18863_ _18863_/A VGND VGND VPWR VPWR _18863_/Y sky130_fd_sc_hd__inv_2
X_17814_ _17914_/A _17812_/X _17814_/C VGND VGND VPWR VPWR _17815_/C sky130_fd_sc_hd__and3_4
X_18794_ _17861_/B VGND VGND VPWR VPWR _18794_/Y sky130_fd_sc_hd__inv_2
X_17745_ _17861_/A _17745_/B VGND VGND VPWR VPWR _17746_/C sky130_fd_sc_hd__or2_4
XFILLER_130_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14957_ _15197_/A _24259_/Q _24678_/Q _14956_/Y VGND VGND VPWR VPWR _14957_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22193__B1 _25199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11563__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13908_ _13908_/A VGND VGND VPWR VPWR _13908_/X sky130_fd_sc_hd__buf_2
XANTENNA__23737__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17676_ _17918_/A VGND VGND VPWR VPWR _17676_/X sky130_fd_sc_hd__buf_2
X_14888_ _24677_/Q VGND VGND VPWR VPWR _14888_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_15_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_30_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19415_ _13032_/B VGND VGND VPWR VPWR _19415_/Y sky130_fd_sc_hd__inv_2
X_16627_ _16627_/A VGND VGND VPWR VPWR _16628_/A sky130_fd_sc_hd__inv_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13839_ _13852_/A _13866_/B _13838_/Y _13867_/C VGND VGND VPWR VPWR _13839_/X sky130_fd_sc_hd__or4_4
XFILLER_56_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19346_ _19345_/Y _19341_/X _19232_/X _19327_/Y VGND VGND VPWR VPWR _19346_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21892__A1_N _14230_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21299__A2 _24257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16558_ _13644_/A VGND VGND VPWR VPWR _16558_/X sky130_fd_sc_hd__buf_2
XFILLER_31_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15509_ _15470_/Y VGND VGND VPWR VPWR _15509_/X sky130_fd_sc_hd__buf_2
X_19277_ _19276_/Y VGND VGND VPWR VPWR _21251_/A sky130_fd_sc_hd__buf_2
XFILLER_91_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16489_ _22883_/A _16486_/X _16246_/X _16486_/X VGND VGND VPWR VPWR _16489_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18228_ _18559_/B VGND VGND VPWR VPWR _18228_/X sky130_fd_sc_hd__buf_2
XFILLER_117_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24596__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18159_ _18159_/A VGND VGND VPWR VPWR _18327_/A sky130_fd_sc_hd__inv_2
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24525__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21170_ _21352_/A _19298_/Y VGND VGND VPWR VPWR _21171_/C sky130_fd_sc_hd__or2_4
Xclkbuf_8_225_0_HCLK clkbuf_8_225_0_HCLK/A VGND VGND VPWR VPWR _24049_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_132_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20121_ _17982_/A _20119_/X _13668_/A _21795_/A _20117_/X VGND VGND VPWR VPWR _23083_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_98_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20052_ _23110_/Q VGND VGND VPWR VPWR _20983_/B sky130_fd_sc_hd__inv_2
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24860_ _23657_/CLK _14085_/X HRESETn VGND VGND VPWR VPWR _14083_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_6_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23811_ _23624_/CLK _18625_/X HRESETn VGND VGND VPWR VPWR _23811_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_96_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24791_ _24823_/CLK _14289_/X HRESETn VGND VGND VPWR VPWR _14286_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12569__A _24510_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23742_ _24182_/CLK _23742_/D HRESETn VGND VGND VPWR VPWR _23742_/Q sky130_fd_sc_hd__dfrtp_4
X_20954_ _18047_/Y VGND VGND VPWR VPWR _22105_/A sky130_fd_sc_hd__buf_2
XANTENNA__20734__A1 sda_oen_o_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23673_ _23680_/CLK _20376_/Y HRESETn VGND VGND VPWR VPWR _20372_/A sky130_fd_sc_hd__dfrtp_4
X_20885_ _12062_/A VGND VGND VPWR VPWR _20885_/X sky130_fd_sc_hd__buf_2
XPHY_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15610__B1 _11573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22624_ _22624_/A _22587_/B VGND VGND VPWR VPWR _22624_/X sky130_fd_sc_hd__and2_4
XPHY_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22555_ _11961_/X VGND VGND VPWR VPWR _22956_/B sky130_fd_sc_hd__buf_2
XANTENNA__21113__C _21113_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21506_ _21211_/A _21506_/B VGND VGND VPWR VPWR _21506_/X sky130_fd_sc_hd__or2_4
X_22486_ _22354_/A _22486_/B VGND VGND VPWR VPWR _22486_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__12304__A2_N _24478_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_35_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_71_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24225_ _24225_/CLK _24225_/D HRESETn VGND VGND VPWR VPWR _16381_/A sky130_fd_sc_hd__dfrtp_4
X_21437_ _24128_/Q _20931_/X _21300_/Y _21436_/X VGND VGND VPWR VPWR _21437_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24266__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12170_ _12170_/A _12170_/B VGND VGND VPWR VPWR _12193_/A sky130_fd_sc_hd__or2_4
XFILLER_120_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24156_ _24104_/CLK _16567_/X HRESETn VGND VGND VPWR VPWR _24156_/Q sky130_fd_sc_hd__dfrtp_4
X_21368_ _21235_/A _19002_/Y VGND VGND VPWR VPWR _21368_/X sky130_fd_sc_hd__or2_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20670__B1 _20647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23107_ _23109_/CLK _20061_/X VGND VGND VPWR VPWR _21649_/C sky130_fd_sc_hd__dfxtp_4
X_20319_ _18617_/X _20318_/Y _20315_/C VGND VGND VPWR VPWR _20319_/X sky130_fd_sc_hd__and3_4
XFILLER_27_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24087_ _24623_/CLK _24087_/D HRESETn VGND VGND VPWR VPWR _16798_/A sky130_fd_sc_hd__dfrtp_4
X_21299_ _21300_/A _24257_/Q _13613_/A VGND VGND VPWR VPWR _21299_/X sky130_fd_sc_hd__o21a_4
XFILLER_1_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23038_ _18005_/Y _21807_/B VGND VGND VPWR VPWR _23038_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__19547__A2_N _19546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15860_ _15847_/A VGND VGND VPWR VPWR _15860_/X sky130_fd_sc_hd__buf_2
XFILLER_40_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14811_ _14806_/X _14807_/X _14808_/X _14811_/D VGND VGND VPWR VPWR _14811_/X sky130_fd_sc_hd__or4_4
X_15791_ _15767_/X VGND VGND VPWR VPWR _15791_/X sky130_fd_sc_hd__buf_2
XANTENNA__12479__A _12412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24989_ _24953_/CLK _24989_/D HRESETn VGND VGND VPWR VPWR _13350_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18918__B2 _18899_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17530_ _17528_/X _17524_/Y _17529_/X VGND VGND VPWR VPWR _17531_/A sky130_fd_sc_hd__or3_4
XANTENNA__23830__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11954_ _11954_/A VGND VGND VPWR VPWR _11954_/X sky130_fd_sc_hd__buf_2
X_14742_ _24691_/Q VGND VGND VPWR VPWR _14742_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25054__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14673_ _24719_/Q _14610_/B _24719_/Q _14610_/B VGND VGND VPWR VPWR _14673_/X sky130_fd_sc_hd__a2bb2o_4
X_17461_ _17453_/X _17460_/X VGND VGND VPWR VPWR _17461_/X sky130_fd_sc_hd__or2_4
X_11885_ _11884_/X VGND VGND VPWR VPWR _11885_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19200_ _17855_/B VGND VGND VPWR VPWR _19200_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15601__B1 _24525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13624_ _13609_/X VGND VGND VPWR VPWR _13624_/Y sky130_fd_sc_hd__inv_2
X_16412_ _16411_/Y _16409_/X _15479_/X _16409_/X VGND VGND VPWR VPWR _24215_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21076__A2_N _20863_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22478__A1 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_117_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_235_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17392_ _17390_/A _17386_/B _17392_/C VGND VGND VPWR VPWR _17392_/X sky130_fd_sc_hd__and3_4
XANTENNA__22478__B2 _22228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19131_ _19129_/Y _19125_/X _19041_/X _19130_/X VGND VGND VPWR VPWR _23444_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20489__B1 _24599_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13555_ _11687_/Y _13555_/B VGND VGND VPWR VPWR _13555_/X sky130_fd_sc_hd__or2_4
X_16343_ _24239_/Q VGND VGND VPWR VPWR _16343_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12506_ _12508_/B VGND VGND VPWR VPWR _12507_/B sky130_fd_sc_hd__inv_2
XANTENNA__13103__A _11741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16274_ _16268_/X _16269_/X _16093_/A _22399_/A _16270_/X VGND VGND VPWR VPWR _16274_/X
+ sky130_fd_sc_hd__a32o_4
X_19062_ _19061_/Y _19058_/X _19038_/X _19058_/X VGND VGND VPWR VPWR _19062_/X sky130_fd_sc_hd__a2bb2o_4
X_13486_ _13468_/A VGND VGND VPWR VPWR _13486_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15225_ _15224_/A _15224_/B VGND VGND VPWR VPWR _15225_/X sky130_fd_sc_hd__or2_4
X_18013_ _23906_/Q VGND VGND VPWR VPWR _18013_/Y sky130_fd_sc_hd__inv_2
X_12437_ _12418_/C _12417_/B VGND VGND VPWR VPWR _12438_/A sky130_fd_sc_hd__or2_4
XFILLER_126_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16414__A _16426_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15156_ _15144_/A _15156_/B _15156_/C VGND VGND VPWR VPWR _15156_/X sky130_fd_sc_hd__or3_4
X_12368_ _12498_/A _24480_/Q _12498_/A _24480_/Q VGND VGND VPWR VPWR _12368_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21453__A2 _11514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15668__B1 _15332_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14107_ _14107_/A VGND VGND VPWR VPWR _14107_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11558__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15087_ _15087_/A _15093_/B VGND VGND VPWR VPWR _15087_/X sky130_fd_sc_hd__or2_4
X_19964_ _19962_/Y _19960_/X _19963_/X _19960_/X VGND VGND VPWR VPWR _23144_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12299_ _12299_/A _12299_/B VGND VGND VPWR VPWR _12300_/B sky130_fd_sc_hd__or2_4
XFILLER_99_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14038_ _14036_/Y _14037_/X _13638_/X _14028_/X VGND VGND VPWR VPWR _24875_/D sky130_fd_sc_hd__a2bb2o_4
X_18915_ _18915_/A VGND VGND VPWR VPWR _18915_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22402__B2 _16305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23989__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19895_ _21513_/B _19890_/X _19828_/X _19890_/X VGND VGND VPWR VPWR _19895_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_55_0_HCLK clkbuf_8_55_0_HCLK/A VGND VGND VPWR VPWR _23949_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_95_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18846_ _21375_/B _18845_/X _15563_/X _18845_/X VGND VGND VPWR VPWR _23545_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23806__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23918__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18777_ _18775_/Y _18776_/X _18706_/X _18776_/X VGND VGND VPWR VPWR _23569_/D sky130_fd_sc_hd__a2bb2o_4
X_15989_ _24365_/Q VGND VGND VPWR VPWR _15989_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22166__B1 _20782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15840__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17728_ _17816_/A _23437_/Q VGND VGND VPWR VPWR _17731_/B sky130_fd_sc_hd__or2_4
XFILLER_36_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20716__A1 sda_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17659_ _17653_/Y _13407_/B _17656_/Y _13407_/A _17658_/X VGND VGND VPWR VPWR _17659_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20670_ _22883_/A _20552_/X _20647_/A _20669_/Y VGND VGND VPWR VPWR _20671_/A sky130_fd_sc_hd__o22a_4
XANTENNA__24777__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19329_ _18763_/X VGND VGND VPWR VPWR _19329_/X sky130_fd_sc_hd__buf_2
XFILLER_108_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24706__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22340_ _24137_/Q _15692_/A _11532_/A _22339_/X VGND VGND VPWR VPWR _22341_/C sky130_fd_sc_hd__a211o_4
XFILLER_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22271_ _22271_/A _20911_/X VGND VGND VPWR VPWR _22271_/X sky130_fd_sc_hd__and2_4
XFILLER_117_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19098__B1 _18964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24010_ _23925_/CLK _17235_/Y HRESETn VGND VGND VPWR VPWR _11728_/C sky130_fd_sc_hd__dfrtp_4
X_21222_ _21234_/A VGND VGND VPWR VPWR _21383_/A sky130_fd_sc_hd__buf_2
XANTENNA__16043__B _23763_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21153_ _21153_/A VGND VGND VPWR VPWR _21159_/A sky130_fd_sc_hd__buf_2
XFILLER_132_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22528__A1_N _12474_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20104_ _20102_/Y _20098_/X _19603_/A _20103_/X VGND VGND VPWR VPWR _20104_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21084_ _20806_/A VGND VGND VPWR VPWR _21425_/B sky130_fd_sc_hd__buf_2
XFILLER_8_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20035_ _20035_/A VGND VGND VPWR VPWR _20035_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23659__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24912_ _24904_/CLK _24912_/D HRESETn VGND VGND VPWR VPWR _13869_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24843_ _24962_/CLK _24843_/D HRESETn VGND VGND VPWR VPWR _24843_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_39_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15831__B1 _11522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24774_ _24776_/CLK _14343_/X HRESETn VGND VGND VPWR VPWR _24774_/Q sky130_fd_sc_hd__dfrtp_4
X_21986_ _22197_/A VGND VGND VPWR VPWR _21986_/X sky130_fd_sc_hd__buf_2
XPHY_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23725_ _24185_/CLK _20548_/X HRESETn VGND VGND VPWR VPWR _20545_/A sky130_fd_sc_hd__dfrtp_4
X_20937_ _16555_/Y _20900_/A VGND VGND VPWR VPWR _20937_/X sky130_fd_sc_hd__and2_4
XPHY_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11670_/A VGND VGND VPWR VPWR _13558_/A sky130_fd_sc_hd__inv_2
XFILLER_39_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21124__B _21590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23656_ _24879_/CLK _20210_/X HRESETn VGND VGND VPWR VPWR _23656_/Q sky130_fd_sc_hd__dfrtp_4
X_20868_ _22444_/B _20858_/X _20864_/Y _20866_/X _20867_/X VGND VGND VPWR VPWR _20868_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_30_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22607_ _12412_/A _22606_/X _24045_/Q _22121_/X VGND VGND VPWR VPWR _22612_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16139__B2 _16138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23587_ _23586_/CLK _18722_/X VGND VGND VPWR VPWR _18721_/A sky130_fd_sc_hd__dfxtp_4
X_20799_ _22148_/A VGND VGND VPWR VPWR _20799_/X sky130_fd_sc_hd__buf_2
XPHY_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24447__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13340_ _13332_/Y _13339_/X _11612_/X _13339_/X VGND VGND VPWR VPWR _24994_/D sky130_fd_sc_hd__a2bb2o_4
X_22538_ _11572_/Y _22536_/X _15957_/Y _22537_/X VGND VGND VPWR VPWR _22538_/X sky130_fd_sc_hd__o22a_4
XFILLER_127_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15898__B1 _15897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21140__A _21144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13271_ _13271_/A _13271_/B _13271_/C VGND VGND VPWR VPWR _13272_/C sky130_fd_sc_hd__or3_4
X_22469_ _24482_/Q _21710_/B VGND VGND VPWR VPWR _22469_/X sky130_fd_sc_hd__or2_4
X_15010_ _14868_/B _15014_/B _14984_/X _15006_/Y VGND VGND VPWR VPWR _15011_/A sky130_fd_sc_hd__a211o_4
X_12222_ _25125_/Q _12222_/B VGND VGND VPWR VPWR _12222_/X sky130_fd_sc_hd__or2_4
X_24208_ _24654_/CLK _16429_/X HRESETn VGND VGND VPWR VPWR _24208_/Q sky130_fd_sc_hd__dfrtp_4
X_25188_ _23353_/CLK _25188_/D HRESETn VGND VGND VPWR VPWR _11698_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12153_ _12152_/Y _24548_/Q _12299_/A _12124_/Y VGND VGND VPWR VPWR _12153_/X sky130_fd_sc_hd__a2bb2o_4
X_24139_ _24113_/CLK _16598_/X HRESETn VGND VGND VPWR VPWR _24139_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12084_ _12083_/X _24561_/Q _12083_/A _24561_/Q VGND VGND VPWR VPWR _12084_/X sky130_fd_sc_hd__a2bb2o_4
X_16961_ _16961_/A VGND VGND VPWR VPWR _17034_/C sky130_fd_sc_hd__inv_2
XFILLER_123_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18700_ _16545_/X VGND VGND VPWR VPWR _18700_/X sky130_fd_sc_hd__buf_2
X_15912_ _15431_/X VGND VGND VPWR VPWR _15912_/X sky130_fd_sc_hd__buf_2
X_19680_ _19680_/A VGND VGND VPWR VPWR _19680_/X sky130_fd_sc_hd__buf_2
XFILLER_103_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16892_ _16891_/X VGND VGND VPWR VPWR _16892_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18631_ _23693_/Q _14349_/Y _20715_/A _20271_/A VGND VGND VPWR VPWR _23805_/D sky130_fd_sc_hd__o22a_4
X_15843_ _15841_/Y _15842_/X _11545_/X _15842_/X VGND VGND VPWR VPWR _15843_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18562_ _16341_/Y _23831_/Q _16341_/Y _23831_/Q VGND VGND VPWR VPWR _18562_/X sky130_fd_sc_hd__a2bb2o_4
X_12986_ _12815_/Y _12984_/X _12985_/Y VGND VGND VPWR VPWR _12986_/X sky130_fd_sc_hd__o21a_4
X_15774_ _12810_/Y _15768_/X _15772_/X _15773_/X VGND VGND VPWR VPWR _15774_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17513_ _17478_/Y _17512_/X _16748_/X _17508_/B VGND VGND VPWR VPWR _17513_/X sky130_fd_sc_hd__a211o_4
X_14725_ _14872_/B VGND VGND VPWR VPWR _15067_/B sky130_fd_sc_hd__buf_2
X_11937_ _11723_/X VGND VGND VPWR VPWR _21300_/B sky130_fd_sc_hd__buf_2
X_18493_ _18488_/A _18488_/B _18475_/X _18489_/Y VGND VGND VPWR VPWR _18494_/A sky130_fd_sc_hd__a211o_4
XANTENNA__16409__A _16426_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17444_ _17323_/D _17366_/X _17345_/X _17441_/Y VGND VGND VPWR VPWR _17445_/A sky130_fd_sc_hd__a211o_4
X_11868_ _11868_/A VGND VGND VPWR VPWR _11868_/Y sky130_fd_sc_hd__inv_2
X_14656_ _14636_/X _14654_/Y _24725_/Q _14655_/X VGND VGND VPWR VPWR _14656_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13607_ _24946_/Q VGND VGND VPWR VPWR _14403_/A sky130_fd_sc_hd__inv_2
X_17375_ _17246_/A _17375_/B VGND VGND VPWR VPWR _17377_/B sky130_fd_sc_hd__or2_4
X_11799_ _11796_/B VGND VGND VPWR VPWR _11799_/Y sky130_fd_sc_hd__inv_2
X_14587_ _14587_/A _19946_/A VGND VGND VPWR VPWR _14587_/X sky130_fd_sc_hd__or2_4
X_19114_ _19114_/A VGND VGND VPWR VPWR _19114_/X sky130_fd_sc_hd__buf_2
XANTENNA__24188__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16326_ _16339_/A VGND VGND VPWR VPWR _16326_/X sky130_fd_sc_hd__buf_2
X_13538_ _13537_/X VGND VGND VPWR VPWR _20660_/B sky130_fd_sc_hd__buf_2
XANTENNA__22871__A1 _21864_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22146__A _14726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12383__A1_N _12416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24117__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19045_ _19044_/Y _19042_/X _18953_/X _19042_/X VGND VGND VPWR VPWR _19045_/X sky130_fd_sc_hd__a2bb2o_4
X_13469_ _13465_/Y _13480_/A _13468_/Y VGND VGND VPWR VPWR _13470_/B sky130_fd_sc_hd__o21ai_4
X_16257_ _16262_/A VGND VGND VPWR VPWR _16257_/X sky130_fd_sc_hd__buf_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15208_ _15208_/A _15211_/B VGND VGND VPWR VPWR _15208_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__21985__A _16202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16188_ _16188_/A VGND VGND VPWR VPWR _16188_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15139_ _15139_/A VGND VGND VPWR VPWR _15144_/B sky130_fd_sc_hd__inv_2
XANTENNA__19455__A _19455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16069__A1_N _16068_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19947_ _19946_/X VGND VGND VPWR VPWR _19960_/A sky130_fd_sc_hd__inv_2
XANTENNA__22926__A2 _15919_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23752__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19878_ _23176_/Q VGND VGND VPWR VPWR _19878_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18829_ _18827_/Y _18822_/X _18828_/X _18809_/A VGND VGND VPWR VPWR _18829_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14749__D _14748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21840_ _21840_/A _15578_/B VGND VGND VPWR VPWR _21840_/X sky130_fd_sc_hd__or2_4
XANTENNA__13008__A _12925_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14962__A2_N _14960_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24958__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21771_ _21519_/A _21769_/X _21771_/C VGND VGND VPWR VPWR _21771_/X sky130_fd_sc_hd__and3_4
XFILLER_36_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21362__B2 _21357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23510_ _23514_/CLK _23510_/D VGND VGND VPWR VPWR _17685_/B sky130_fd_sc_hd__dfxtp_4
X_20722_ _14633_/X _20721_/X _20729_/B VGND VGND VPWR VPWR _23686_/D sky130_fd_sc_hd__o21a_4
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24490_ _24307_/CLK _15675_/X HRESETn VGND VGND VPWR VPWR _24490_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23441_ _23479_/CLK _19138_/X VGND VGND VPWR VPWR _19136_/A sky130_fd_sc_hd__dfxtp_4
X_20653_ _20653_/A _20653_/B VGND VGND VPWR VPWR _20653_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__13052__B1 _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_100_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_201_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24540__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11602__A1 _11533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23372_ _23374_/CLK _19335_/X VGND VGND VPWR VPWR _19333_/A sky130_fd_sc_hd__dfxtp_4
X_20584_ _13533_/A VGND VGND VPWR VPWR _20584_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25111_ _25115_/CLK _12278_/X HRESETn VGND VGND VPWR VPWR _12110_/A sky130_fd_sc_hd__dfrtp_4
X_22323_ _22323_/A _22188_/X VGND VGND VPWR VPWR _22323_/X sky130_fd_sc_hd__and2_4
XFILLER_30_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12582__A _12582_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16054__A _16054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25042_ _25044_/CLK _12759_/X HRESETn VGND VGND VPWR VPWR _12593_/A sky130_fd_sc_hd__dfrtp_4
X_22254_ _22919_/A _22242_/X _22245_/X _22254_/D VGND VGND VPWR VPWR _22254_/X sky130_fd_sc_hd__or4_4
XANTENNA__18818__B1 _18817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21205_ _21205_/A VGND VGND VPWR VPWR _21371_/A sky130_fd_sc_hd__buf_2
XANTENNA__20625__B1 _24173_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21968__A3 _21938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22185_ _22155_/A _22184_/X _21046_/X _24554_/Q _22884_/B VGND VGND VPWR VPWR _22185_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21136_ _17651_/A VGND VGND VPWR VPWR _21469_/A sky130_fd_sc_hd__buf_2
XFILLER_120_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22378__B1 _24039_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15831__A1_N _15830_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21067_ _13499_/A VGND VGND VPWR VPWR _21067_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16057__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20018_ _21917_/B _20015_/X _19714_/X _20015_/X VGND VGND VPWR VPWR _20018_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14021__B _20852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12840_ _12951_/A VGND VGND VPWR VPWR _12947_/A sky130_fd_sc_hd__inv_2
XFILLER_104_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24826_ _24824_/CLK _24826_/D HRESETn VGND VGND VPWR VPWR _24826_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24699__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12771_ _12762_/X _12770_/X _12755_/X VGND VGND VPWR VPWR _25038_/D sky130_fd_sc_hd__and3_4
X_21969_ _21062_/X _21968_/X VGND VGND VPWR VPWR _22004_/C sky130_fd_sc_hd__nor2_4
XANTENNA__18143__A1_N _24345_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24757_ _24757_/CLK _14418_/X HRESETn VGND VGND VPWR VPWR _14377_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22550__B1 _14933_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11499_/A VGND VGND VPWR VPWR _13612_/A sky130_fd_sc_hd__inv_2
X_14510_ _14509_/X VGND VGND VPWR VPWR _14510_/Y sky130_fd_sc_hd__inv_2
XPHY_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15472_/A VGND VGND VPWR VPWR _15490_/X sky130_fd_sc_hd__buf_2
X_23708_ _23706_/CLK _23708_/D HRESETn VGND VGND VPWR VPWR _13508_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_15_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24688_ _24712_/CLK _24688_/D HRESETn VGND VGND VPWR VPWR _24688_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20974__A _20979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11653_/A VGND VGND VPWR VPWR _13571_/A sky130_fd_sc_hd__inv_2
X_14441_ _14441_/A VGND VGND VPWR VPWR _21012_/A sky130_fd_sc_hd__buf_2
XFILLER_39_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23639_ _24811_/CLK _20321_/Y HRESETn VGND VGND VPWR VPWR _18617_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_42_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21105__B2 _21050_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24281__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14372_ _14372_/A VGND VGND VPWR VPWR _14387_/A sky130_fd_sc_hd__buf_2
X_17160_ _17160_/A _17160_/B VGND VGND VPWR VPWR _17161_/B sky130_fd_sc_hd__or2_4
XPHY_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11584_ HWDATA[14] VGND VGND VPWR VPWR _11585_/A sky130_fd_sc_hd__buf_2
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19259__B _23763_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24210__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13323_ _24619_/Q VGND VGND VPWR VPWR _14195_/B sky130_fd_sc_hd__buf_2
X_16111_ _16111_/A VGND VGND VPWR VPWR _21858_/A sky130_fd_sc_hd__inv_2
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17091_ _17044_/X _17054_/B _17076_/A VGND VGND VPWR VPWR _17092_/C sky130_fd_sc_hd__o21a_4
XFILLER_122_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13254_ _13222_/A _13250_/X _13254_/C VGND VGND VPWR VPWR _13254_/X sky130_fd_sc_hd__or3_4
X_16042_ _16042_/A VGND VGND VPWR VPWR _22265_/B sky130_fd_sc_hd__buf_2
XFILLER_136_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12205_ _12204_/X VGND VGND VPWR VPWR _12205_/Y sky130_fd_sc_hd__inv_2
X_13185_ _11751_/X VGND VGND VPWR VPWR _13221_/A sky130_fd_sc_hd__buf_2
X_19801_ _19801_/A _19801_/B VGND VGND VPWR VPWR _19802_/A sky130_fd_sc_hd__nand2_4
XFILLER_69_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12136_ _25119_/Q VGND VGND VPWR VPWR _12174_/B sky130_fd_sc_hd__inv_2
X_17993_ HWDATA[7] VGND VGND VPWR VPWR _17993_/X sky130_fd_sc_hd__buf_2
XFILLER_97_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19732_ _21132_/B _19727_/X _19731_/X _19727_/X VGND VGND VPWR VPWR _19732_/X sky130_fd_sc_hd__a2bb2o_4
X_12067_ _11956_/X _16302_/A VGND VGND VPWR VPWR _12067_/Y sky130_fd_sc_hd__nor2_4
X_16944_ _16924_/B _16943_/X _16951_/C VGND VGND VPWR VPWR _24064_/D sky130_fd_sc_hd__and3_4
X_19663_ _19663_/A VGND VGND VPWR VPWR _20984_/B sky130_fd_sc_hd__inv_2
X_16875_ _16867_/A _16875_/B _16874_/Y VGND VGND VPWR VPWR _16875_/X sky130_fd_sc_hd__and3_4
XFILLER_38_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12135__A2_N _24568_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18614_ _18614_/A _18614_/B VGND VGND VPWR VPWR _18614_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_129_0_HCLK clkbuf_7_64_0_HCLK/X VGND VGND VPWR VPWR _23457_/CLK sky130_fd_sc_hd__clkbuf_1
X_15826_ _15826_/A VGND VGND VPWR VPWR _15826_/X sky130_fd_sc_hd__buf_2
X_19594_ _23278_/Q VGND VGND VPWR VPWR _19594_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21045__A _21034_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19537__B2 _19534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18545_ _18545_/A VGND VGND VPWR VPWR _18546_/B sky130_fd_sc_hd__inv_2
X_15757_ _15757_/A VGND VGND VPWR VPWR _15757_/X sky130_fd_sc_hd__buf_2
X_12969_ _12964_/A _12964_/B _12922_/X _12965_/Y VGND VGND VPWR VPWR _12969_/X sky130_fd_sc_hd__a211o_4
XFILLER_45_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24369__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14708_ _15033_/A _22502_/A _14876_/D _22502_/A VGND VGND VPWR VPWR _14708_/X sky130_fd_sc_hd__a2bb2o_4
X_18476_ _18470_/A _18470_/B _18475_/X _18472_/B VGND VGND VPWR VPWR _18476_/X sky130_fd_sc_hd__a211o_4
X_15688_ _15684_/X _15672_/X _15499_/X _24481_/Q _15685_/X VGND VGND VPWR VPWR _15688_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16220__B1 _16219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17427_ _17300_/X VGND VGND VPWR VPWR _17428_/C sky130_fd_sc_hd__buf_2
XANTENNA__15978__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14639_ _14639_/A VGND VGND VPWR VPWR _14639_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17358_ _17255_/Y _17358_/B VGND VGND VPWR VPWR _17362_/B sky130_fd_sc_hd__or2_4
X_16309_ _16304_/Y _16308_/X _15828_/X _16308_/X VGND VGND VPWR VPWR _24253_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17289_ _25212_/Q _17288_/Y _11562_/Y _23998_/Q VGND VGND VPWR VPWR _17289_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19028_ _21209_/B _19025_/X _15566_/X _19025_/X VGND VGND VPWR VPWR _19028_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19301__A2_N _19296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23933__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25157__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16287__B1 _15897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22323__B _22188_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14837__B2 _14836_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23990_ _23990_/CLK _17406_/Y HRESETn VGND VGND VPWR VPWR _23990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_25_0_HCLK clkbuf_6_12_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22941_ _12579_/Y _20910_/X _12813_/Y _22029_/X VGND VGND VPWR VPWR _22941_/X sky130_fd_sc_hd__o22a_4
XFILLER_25_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14271__A2_N _14268_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_88_0_HCLK clkbuf_6_44_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_88_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__22780__B1 _20801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20778__B _20777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22872_ _13337_/A _22868_/Y _22407_/X _22871_/X VGND VGND VPWR VPWR _22872_/X sky130_fd_sc_hd__o22a_4
XFILLER_84_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21823_ _20965_/A VGND VGND VPWR VPWR _21913_/A sky130_fd_sc_hd__buf_2
XFILLER_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24792__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24611_ _24182_/CLK _24611_/D HRESETn VGND VGND VPWR VPWR _24611_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22993__B _22870_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24721__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24542_ _24618_/CLK _15532_/X HRESETn VGND VGND VPWR VPWR _13519_/A sky130_fd_sc_hd__dfrtp_4
X_21754_ _21753_/X VGND VGND VPWR VPWR _21754_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20794__A _22501_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24039__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20705_ _23808_/Q _20705_/B VGND VGND VPWR VPWR _20705_/X sky130_fd_sc_hd__and2_4
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24473_ _24307_/CLK _15701_/X HRESETn VGND VGND VPWR VPWR _24473_/Q sky130_fd_sc_hd__dfrtp_4
X_21685_ _22064_/A _19824_/Y VGND VGND VPWR VPWR _21685_/X sky130_fd_sc_hd__or2_4
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23424_ _23425_/CLK _23424_/D VGND VGND VPWR VPWR _23424_/Q sky130_fd_sc_hd__dfxtp_4
X_20636_ _20634_/Y _20631_/X _20635_/X VGND VGND VPWR VPWR _20636_/X sky130_fd_sc_hd__o21a_4
XFILLER_138_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23355_ _23350_/CLK _19382_/X VGND VGND VPWR VPWR _19380_/A sky130_fd_sc_hd__dfxtp_4
X_20567_ _20566_/Y _13528_/A _13529_/X VGND VGND VPWR VPWR _20567_/X sky130_fd_sc_hd__o21a_4
X_22306_ _22306_/A _22296_/X _22299_/X _22305_/X VGND VGND VPWR VPWR _22306_/X sky130_fd_sc_hd__or4_4
X_23286_ _23308_/CLK _19577_/X VGND VGND VPWR VPWR _19573_/A sky130_fd_sc_hd__dfxtp_4
X_20498_ _20499_/B VGND VGND VPWR VPWR _20498_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22514__A _21848_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25025_ _25021_/CLK _25025_/D HRESETn VGND VGND VPWR VPWR _12854_/A sky130_fd_sc_hd__dfrtp_4
X_22237_ _21642_/X VGND VGND VPWR VPWR _22919_/A sky130_fd_sc_hd__buf_2
XFILLER_3_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23674__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22168_ _22168_/A _22163_/X _22168_/C VGND VGND VPWR VPWR _22168_/X sky130_fd_sc_hd__or3_4
XANTENNA__14828__A1 _24695_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21119_ _11952_/X _21118_/X VGND VGND VPWR VPWR _21119_/X sky130_fd_sc_hd__or2_4
XANTENNA__19216__B1 _19149_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14990_ _14990_/A _14990_/B VGND VGND VPWR VPWR _14991_/C sky130_fd_sc_hd__or2_4
X_22099_ _20964_/A _19686_/Y VGND VGND VPWR VPWR _22101_/B sky130_fd_sc_hd__or2_4
XFILLER_120_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21023__B1 _13334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13941_ _13926_/C _13941_/B _13927_/A VGND VGND VPWR VPWR _13941_/X sky130_fd_sc_hd__or3_4
XFILLER_130_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21574__A1 _24129_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16660_ _16658_/Y _16650_/X _15507_/X _16659_/X VGND VGND VPWR VPWR _16660_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13872_ _13872_/A _13871_/X _13872_/C _13851_/B VGND VGND VPWR VPWR _13873_/A sky130_fd_sc_hd__or4_4
XFILLER_62_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18082__A1_N _13011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15611_ _16624_/A VGND VGND VPWR VPWR _15611_/X sky130_fd_sc_hd__buf_2
X_12823_ _24446_/Q VGND VGND VPWR VPWR _12823_/Y sky130_fd_sc_hd__inv_2
X_24809_ _24788_/CLK _14245_/X HRESETn VGND VGND VPWR VPWR _24809_/Q sky130_fd_sc_hd__dfstp_4
X_16591_ _16581_/X _16573_/X HWDATA[18] _24143_/Q _16590_/X VGND VGND VPWR VPWR _16591_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_76_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18330_ _18328_/Y _18329_/X _18319_/X VGND VGND VPWR VPWR _23848_/D sky130_fd_sc_hd__and3_4
XANTENNA__24462__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15542_ _15540_/Y _15537_/X _15541_/X _15537_/X VGND VGND VPWR VPWR _24540_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12754_ _12739_/A _12739_/B VGND VGND VPWR VPWR _12754_/Y sky130_fd_sc_hd__nand2_4
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21877__A2 _21082_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11705_ _11698_/C VGND VGND VPWR VPWR _18638_/A sky130_fd_sc_hd__inv_2
X_18261_ _18260_/X VGND VGND VPWR VPWR _23867_/D sky130_fd_sc_hd__inv_2
XPHY_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _13007_/B _12685_/B _12685_/C VGND VGND VPWR VPWR _12686_/A sky130_fd_sc_hd__or3_4
X_15473_ _12108_/Y _15472_/X _11525_/X _15472_/X VGND VGND VPWR VPWR _15473_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _24014_/Q VGND VGND VPWR VPWR _17212_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22408__B _22188_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ _15801_/A VGND VGND VPWR VPWR _11636_/X sky130_fd_sc_hd__buf_2
X_14424_ _14424_/A _14424_/B VGND VGND VPWR VPWR _14424_/X sky130_fd_sc_hd__or2_4
XANTENNA__14764__B1 _15019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18192_ _18164_/X _18192_/B VGND VGND VPWR VPWR _18485_/C sky130_fd_sc_hd__or2_4
XFILLER_30_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11578__B1 _11576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17143_ _17143_/A VGND VGND VPWR VPWR _17143_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14807__A2_N _24125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11567_ _11565_/Y _11559_/X _11566_/X _11559_/X VGND VGND VPWR VPWR _25209_/D sky130_fd_sc_hd__a2bb2o_4
X_14355_ _20185_/A _14355_/B VGND VGND VPWR VPWR _24771_/D sky130_fd_sc_hd__or2_4
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13306_ _13085_/A _13306_/B VGND VGND VPWR VPWR _13306_/X sky130_fd_sc_hd__or2_4
X_14286_ _14286_/A VGND VGND VPWR VPWR _14286_/Y sky130_fd_sc_hd__inv_2
X_17074_ _17074_/A _17074_/B _17073_/X VGND VGND VPWR VPWR _17074_/X sky130_fd_sc_hd__or3_4
X_11498_ _24616_/Q VGND VGND VPWR VPWR _12060_/A sky130_fd_sc_hd__inv_2
XANTENNA__22424__A _12362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13237_ _13301_/A _23201_/Q VGND VGND VPWR VPWR _13237_/X sky130_fd_sc_hd__or2_4
X_16025_ _14560_/A _16023_/X _14560_/Y _16024_/Y VGND VGND VPWR VPWR _16027_/A sky130_fd_sc_hd__o22a_4
XFILLER_83_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17518__A _16710_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13168_ _13204_/A _23603_/Q VGND VGND VPWR VPWR _13168_/X sky130_fd_sc_hd__or2_4
XFILLER_83_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12119_ _12119_/A _12119_/B _12115_/X _12118_/X VGND VGND VPWR VPWR _12119_/X sky130_fd_sc_hd__or4_4
XANTENNA__11566__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23003__A1 _22335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15038__A _24699_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13099_ _13316_/A _23381_/Q VGND VGND VPWR VPWR _13099_/X sky130_fd_sc_hd__or2_4
X_17976_ _17975_/Y VGND VGND VPWR VPWR _17987_/A sky130_fd_sc_hd__buf_2
XFILLER_97_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23003__B2 _22576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20879__A _22859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12074__A2_N _24576_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19715_ _21916_/B _19710_/X _19714_/X _19710_/X VGND VGND VPWR VPWR _23237_/D sky130_fd_sc_hd__a2bb2o_4
X_16927_ _16927_/A _16936_/B VGND VGND VPWR VPWR _16927_/X sky130_fd_sc_hd__or2_4
XFILLER_66_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19646_ _19646_/A VGND VGND VPWR VPWR _19646_/Y sky130_fd_sc_hd__inv_2
X_16858_ _16858_/A VGND VGND VPWR VPWR _16858_/X sky130_fd_sc_hd__buf_2
XFILLER_66_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15809_ _15807_/X VGND VGND VPWR VPWR _15810_/B sky130_fd_sc_hd__inv_2
XFILLER_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19577_ _19573_/Y _19576_/X _19442_/X _19576_/X VGND VGND VPWR VPWR _19577_/X sky130_fd_sc_hd__a2bb2o_4
X_16789_ _15877_/Y _24071_/Q _15877_/Y _24071_/Q VGND VGND VPWR VPWR _16789_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18528_ _18338_/X _18527_/Y VGND VGND VPWR VPWR _18530_/B sky130_fd_sc_hd__or2_4
XANTENNA__24132__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18459_ _18459_/A _18438_/X VGND VGND VPWR VPWR _18460_/A sky130_fd_sc_hd__or2_4
XANTENNA__13005__B _13008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15501__A HWDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21470_ _21336_/A _19609_/Y VGND VGND VPWR VPWR _21470_/X sky130_fd_sc_hd__or2_4
XFILLER_18_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20119__A _22218_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20421_ _20420_/X VGND VGND VPWR VPWR _20421_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19240__A2_N _19239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13021__A _13299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23140_ _23332_/CLK _19976_/X VGND VGND VPWR VPWR _23140_/Q sky130_fd_sc_hd__dfxtp_4
X_20352_ _20352_/A VGND VGND VPWR VPWR _20352_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23071_ _23992_/CLK _23071_/D VGND VGND VPWR VPWR _20147_/A sky130_fd_sc_hd__dfxtp_4
X_20283_ _20283_/A _20282_/Y _20278_/X VGND VGND VPWR VPWR _20283_/X sky130_fd_sc_hd__and3_4
XANTENNA__16332__A _24243_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22022_ _22022_/A VGND VGND VPWR VPWR _22022_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22596__A3 _21981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16275__A3 _15505_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24973__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23973_ _24361_/CLK _17509_/X HRESETn VGND VGND VPWR VPWR _23012_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_68_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21556__B2 _20744_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24902__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22924_ _14777_/A _22857_/B VGND VGND VPWR VPWR _22924_/X sky130_fd_sc_hd__or2_4
XFILLER_60_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_112_0_HCLK clkbuf_7_56_0_HCLK/X VGND VGND VPWR VPWR _23657_/CLK sky130_fd_sc_hd__clkbuf_1
X_22855_ _12416_/A _22259_/X _24053_/Q _22433_/A VGND VGND VPWR VPWR _22856_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16983__A1 _24308_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_175_0_HCLK clkbuf_7_87_0_HCLK/X VGND VGND VPWR VPWR _25112_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21806_ _21803_/Y _21804_/X _21649_/X _21805_/X VGND VGND VPWR VPWR _21807_/B sky130_fd_sc_hd__a211o_4
XANTENNA__21859__A2 _21858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22786_ _12448_/A _22259_/A _17026_/B _20747_/X VGND VGND VPWR VPWR _22786_/X sky130_fd_sc_hd__o22a_4
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21737_ _21737_/A _21734_/X _21737_/C _21737_/D VGND VGND VPWR VPWR _21738_/A sky130_fd_sc_hd__or4_4
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24525_ _24483_/CLK _15601_/X HRESETn VGND VGND VPWR VPWR _24525_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22711__A2_N _22708_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15411__A _15410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12470_ _12410_/Y _12468_/A VGND VGND VPWR VPWR _12470_/X sky130_fd_sc_hd__or2_4
X_21668_ _21667_/X _18652_/Y VGND VGND VPWR VPWR _21668_/X sky130_fd_sc_hd__or2_4
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24456_ _24432_/CLK _15758_/X HRESETn VGND VGND VPWR VPWR _22891_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_36_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20619_ _20617_/Y _20614_/Y _20618_/X VGND VGND VPWR VPWR _20619_/X sky130_fd_sc_hd__o21a_4
X_23407_ _23979_/CLK _23407_/D VGND VGND VPWR VPWR _19231_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__23855__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24387_ _24361_/CLK _24387_/D HRESETn VGND VGND VPWR VPWR _24387_/Q sky130_fd_sc_hd__dfrtp_4
X_21599_ _21598_/X VGND VGND VPWR VPWR _21599_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25079__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14140_ _14126_/A _14139_/X _13350_/A _14131_/X VGND VGND VPWR VPWR _24843_/D sky130_fd_sc_hd__o22a_4
X_23338_ _24750_/CLK _23338_/D VGND VGND VPWR VPWR _19429_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__25008__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14071_ _13797_/A _13777_/D _13787_/Y _14071_/D VGND VGND VPWR VPWR _14071_/X sky130_fd_sc_hd__or4_4
XFILLER_10_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15171__B1 _15147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19437__B1 _19392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23269_ _23278_/CLK _23269_/D VGND VGND VPWR VPWR _23269_/Q sky130_fd_sc_hd__dfxtp_4
X_13022_ _13045_/A _13022_/B VGND VGND VPWR VPWR _13022_/X sky130_fd_sc_hd__or2_4
X_25008_ _25009_/CLK _25008_/D HRESETn VGND VGND VPWR VPWR _25008_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_121_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17830_ _17929_/A _17830_/B _17829_/X VGND VGND VPWR VPWR _17830_/X sky130_fd_sc_hd__and3_4
X_17761_ _17903_/A _17761_/B VGND VGND VPWR VPWR _17761_/X sky130_fd_sc_hd__or2_4
X_14973_ _14943_/X _14973_/B _14973_/C _14972_/X VGND VGND VPWR VPWR _14973_/X sky130_fd_sc_hd__or4_4
X_19500_ _23313_/Q VGND VGND VPWR VPWR _19500_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21547__B2 _21544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16712_ _22202_/A VGND VGND VPWR VPWR _16712_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24643__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13924_ _13924_/A VGND VGND VPWR VPWR _13933_/A sky130_fd_sc_hd__inv_2
XFILLER_75_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17692_ _14569_/A _17690_/X _17692_/C VGND VGND VPWR VPWR _17692_/X sky130_fd_sc_hd__and3_4
XFILLER_74_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_71_0_HCLK clkbuf_7_71_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_71_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19431_ _13251_/B VGND VGND VPWR VPWR _19431_/Y sky130_fd_sc_hd__inv_2
X_16643_ _16643_/A VGND VGND VPWR VPWR _16643_/X sky130_fd_sc_hd__buf_2
XFILLER_78_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13855_ _13824_/X _13825_/X _13833_/A VGND VGND VPWR VPWR _13855_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_63_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16974__A1 _16172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13106__A _13309_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12806_ _22126_/A VGND VGND VPWR VPWR _12806_/Y sky130_fd_sc_hd__inv_2
X_19362_ _19362_/A VGND VGND VPWR VPWR _19362_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17801__A _14569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16574_ _15799_/X _16573_/X HWDATA[28] _24153_/Q _16566_/X VGND VGND VPWR VPWR _16574_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_90_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14985__B1 _14984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13786_ _13786_/A VGND VGND VPWR VPWR _13786_/Y sky130_fd_sc_hd__inv_2
X_18313_ _18290_/X _18307_/B _18312_/Y VGND VGND VPWR VPWR _23854_/D sky130_fd_sc_hd__and3_4
X_15525_ _12124_/Y _15518_/X _14304_/X _15472_/A VGND VGND VPWR VPWR _15525_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12737_ _12737_/A _12737_/B VGND VGND VPWR VPWR _12737_/X sky130_fd_sc_hd__or2_4
X_19293_ _23386_/Q VGND VGND VPWR VPWR _19293_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20522__A2 _20416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22138__B _22051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18244_ _18244_/A _18248_/B VGND VGND VPWR VPWR _18246_/B sky130_fd_sc_hd__or2_4
X_15456_ _15455_/X VGND VGND VPWR VPWR _15456_/X sky130_fd_sc_hd__buf_2
X_12668_ _12668_/A VGND VGND VPWR VPWR _25067_/D sky130_fd_sc_hd__inv_2
XANTENNA__11991__A1_N _11985_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ _13438_/Y _14382_/B VGND VGND VPWR VPWR _14407_/Y sky130_fd_sc_hd__nand2_4
X_11619_ HWDATA[5] VGND VGND VPWR VPWR _13668_/A sky130_fd_sc_hd__buf_2
X_18175_ _16080_/Y _23862_/Q _24345_/Q _18268_/A VGND VGND VPWR VPWR _18175_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15387_ _15358_/X VGND VGND VPWR VPWR _15387_/X sky130_fd_sc_hd__buf_2
X_12599_ _12728_/A _24514_/Q _12728_/A _24514_/Q VGND VGND VPWR VPWR _12599_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20881__B _20931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17126_ _17126_/A VGND VGND VPWR VPWR _17127_/B sky130_fd_sc_hd__inv_2
XFILLER_129_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14338_ _21549_/A _14325_/X _21443_/A _14327_/X VGND VGND VPWR VPWR _14338_/X sky130_fd_sc_hd__o22a_4
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17057_ _17056_/Y VGND VGND VPWR VPWR _17057_/X sky130_fd_sc_hd__buf_2
XANTENNA__19428__B1 _19381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14269_ _14266_/X _14268_/X _14228_/X _14268_/X VGND VGND VPWR VPWR _14269_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16152__A _16165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16008_ _14435_/B _15439_/X VGND VGND VPWR VPWR _16008_/X sky130_fd_sc_hd__or2_4
XANTENNA__21993__A _24366_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16662__B1 _16451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17959_ _17927_/A _23455_/Q VGND VGND VPWR VPWR _17959_/X sky130_fd_sc_hd__or2_4
XFILLER_39_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13476__B1 _13480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24384__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20970_ _17642_/Y VGND VGND VPWR VPWR _20975_/A sky130_fd_sc_hd__buf_2
XFILLER_93_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24313__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19629_ _19636_/A VGND VGND VPWR VPWR _19629_/X sky130_fd_sc_hd__buf_2
XFILLER_93_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16965__B2 _17041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13016__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22640_ _22197_/A VGND VGND VPWR VPWR _22640_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_248_0_HCLK clkbuf_7_124_0_HCLK/X VGND VGND VPWR VPWR _24094_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16972__D _16972_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22571_ _22571_/A VGND VGND VPWR VPWR _22572_/C sky130_fd_sc_hd__inv_2
XFILLER_33_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21522_ _21235_/A _21522_/B VGND VGND VPWR VPWR _21522_/X sky130_fd_sc_hd__or2_4
XFILLER_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24310_ _24606_/CLK _24310_/D HRESETn VGND VGND VPWR VPWR _24310_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14256__A1_N _14255_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24241_ _24262_/CLK _24241_/D HRESETn VGND VGND VPWR VPWR _24241_/Q sky130_fd_sc_hd__dfrtp_4
X_21453_ _17487_/Y _11514_/X _12858_/X _15576_/X VGND VGND VPWR VPWR _21453_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21445__A1_N _14257_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25172__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20404_ _23772_/Q _20404_/B _20403_/X VGND VGND VPWR VPWR _20404_/X sky130_fd_sc_hd__and3_4
X_24172_ _24168_/CLK _16521_/X HRESETn VGND VGND VPWR VPWR _16520_/A sky130_fd_sc_hd__dfrtp_4
X_21384_ _21224_/A _21384_/B _21384_/C VGND VGND VPWR VPWR _21384_/X sky130_fd_sc_hd__and3_4
XFILLER_134_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20071__A1_N _21181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25101__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23123_ _23292_/CLK _23123_/D VGND VGND VPWR VPWR _20019_/A sky130_fd_sc_hd__dfxtp_4
X_20335_ _20164_/B VGND VGND VPWR VPWR _20335_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23054_ _23041_/X VGND VGND VPWR VPWR IRQ[2] sky130_fd_sc_hd__buf_2
X_20266_ _20266_/A _20264_/X _20266_/C _20266_/D VGND VGND VPWR VPWR _20266_/X sky130_fd_sc_hd__or4_4
X_22005_ _16457_/Y _22230_/A _14732_/A _21570_/X VGND VGND VPWR VPWR _22005_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19373__A _19372_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20197_ _23761_/D VGND VGND VPWR VPWR _20197_/X sky130_fd_sc_hd__buf_2
XFILLER_88_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21408__A _24470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14824__A1_N _14997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11970_ _25153_/Q VGND VGND VPWR VPWR _11970_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23956_ _23957_/CLK _23956_/D HRESETn VGND VGND VPWR VPWR _22434_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16405__B1 _11536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24054__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_58_0_HCLK clkbuf_6_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_58_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22907_ _24317_/Q _22834_/B VGND VGND VPWR VPWR _22907_/X sky130_fd_sc_hd__or2_4
XANTENNA__15759__A2 _15740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23887_ _25186_/CLK _23887_/D HRESETn VGND VGND VPWR VPWR _21644_/A sky130_fd_sc_hd__dfrtp_4
X_13640_ _13637_/Y _13631_/X _13638_/X _13639_/X VGND VGND VPWR VPWR _24943_/D sky130_fd_sc_hd__a2bb2o_4
X_22838_ _22838_/A _23008_/B VGND VGND VPWR VPWR _22838_/X sky130_fd_sc_hd__or2_4
XFILLER_112_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21143__A _21336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _13571_/A _13564_/X VGND VGND VPWR VPWR _13571_/X sky130_fd_sc_hd__or2_4
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22769_ _22769_/A _22651_/B VGND VGND VPWR VPWR _22769_/X sky130_fd_sc_hd__and2_4
XFILLER_9_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15310_ _15300_/Y VGND VGND VPWR VPWR _15310_/X sky130_fd_sc_hd__buf_2
XFILLER_34_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ _12408_/C _12505_/B VGND VGND VPWR VPWR _12523_/C sky130_fd_sc_hd__nand2_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24508_ _25034_/CLK _15627_/X HRESETn VGND VGND VPWR VPWR _24508_/Q sky130_fd_sc_hd__dfrtp_4
X_16290_ HWDATA[2] VGND VGND VPWR VPWR _16291_/A sky130_fd_sc_hd__buf_2
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19147__A2_N _19146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15241_ _15241_/A VGND VGND VPWR VPWR _15262_/A sky130_fd_sc_hd__inv_2
XFILLER_40_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19777__A2_N _19772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12453_ _12444_/A VGND VGND VPWR VPWR _12453_/X sky130_fd_sc_hd__buf_2
X_24439_ _24502_/CLK _15789_/X HRESETn VGND VGND VPWR VPWR _22243_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18452__A _18459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21465__B1 _18049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12384_ _22736_/A VGND VGND VPWR VPWR _12384_/Y sky130_fd_sc_hd__inv_2
X_15172_ _15105_/A _15170_/X _15171_/Y VGND VGND VPWR VPWR _24669_/D sky130_fd_sc_hd__o21a_4
X_14123_ _14111_/C _14110_/X _13488_/X _14122_/X VGND VGND VPWR VPWR _14124_/A sky130_fd_sc_hd__a211o_4
XFILLER_125_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19980_ _21521_/B _19975_/X _19455_/A _19975_/X VGND VGND VPWR VPWR _19980_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22009__A2 _20819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24627__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14498__A2 _14506_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18931_ _17870_/B VGND VGND VPWR VPWR _18931_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24895__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14054_ _14052_/Y _14048_/X _13668_/X _14053_/X VGND VGND VPWR VPWR _24869_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13005_ _12999_/A _13008_/B VGND VGND VPWR VPWR _13005_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24824__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18862_ _18861_/Y _18859_/X _18817_/X _18859_/X VGND VGND VPWR VPWR _18862_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16239__A3 _15468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17813_ _17881_/A _19955_/A VGND VGND VPWR VPWR _17814_/C sky130_fd_sc_hd__or2_4
XANTENNA__16644__B1 _16261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19715__A2_N _19710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18793_ _18792_/Y _18790_/X _18700_/X _18790_/X VGND VGND VPWR VPWR _23563_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16960__A1_N _16133_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17744_ _17721_/A VGND VGND VPWR VPWR _17861_/A sky130_fd_sc_hd__buf_2
X_14956_ _14956_/A VGND VGND VPWR VPWR _14956_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22193__B2 _22858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13907_ _23691_/Q _13896_/X _13900_/X _24905_/Q _13903_/X VGND VGND VPWR VPWR _13907_/X
+ sky130_fd_sc_hd__a32o_4
X_17675_ _17726_/A VGND VGND VPWR VPWR _17918_/A sky130_fd_sc_hd__buf_2
XANTENNA__12044__A1_N _11985_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14887_ _24261_/Q VGND VGND VPWR VPWR _14887_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19414_ _19413_/Y _19409_/X _19392_/X _19396_/Y VGND VGND VPWR VPWR _23343_/D sky130_fd_sc_hd__a2bb2o_4
X_16626_ _16624_/X _16625_/X HWDATA[30] _24123_/Q _16622_/X VGND VGND VPWR VPWR _16626_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13838_ _13867_/A VGND VGND VPWR VPWR _13838_/Y sky130_fd_sc_hd__inv_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19345_ _13305_/B VGND VGND VPWR VPWR _19345_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21053__A _21590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16557_ _16555_/Y _16493_/A _16556_/X _16493_/A VGND VGND VPWR VPWR _16557_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23777__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_1_0_HCLK clkbuf_6_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_1_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_13769_ _13769_/A _13769_/B _13769_/C _13769_/D VGND VGND VPWR VPWR _13778_/A sky130_fd_sc_hd__or4_4
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_15_0_HCLK clkbuf_7_7_0_HCLK/X VGND VGND VPWR VPWR _23350_/CLK sky130_fd_sc_hd__clkbuf_1
X_15508_ _15503_/X _15504_/X _15507_/X _24556_/Q _15466_/A VGND VGND VPWR VPWR _15508_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_91_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19276_ _23392_/Q VGND VGND VPWR VPWR _19276_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23706__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16488_ _16488_/A VGND VGND VPWR VPWR _22883_/A sky130_fd_sc_hd__inv_2
XANTENNA__20892__A _22018_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_78_0_HCLK clkbuf_8_79_0_HCLK/A VGND VGND VPWR VPWR _23885_/CLK sky130_fd_sc_hd__clkbuf_1
X_18227_ _18262_/A VGND VGND VPWR VPWR _18559_/B sky130_fd_sc_hd__inv_2
XFILLER_31_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15439_ _13454_/X VGND VGND VPWR VPWR _15439_/X sky130_fd_sc_hd__buf_2
XFILLER_50_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15986__A _24366_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20259__A1 _23766_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18158_ _24333_/Q _23854_/Q _22232_/A _18312_/A VGND VGND VPWR VPWR _18158_/X sky130_fd_sc_hd__o22a_4
X_17109_ _17042_/A _17108_/X VGND VGND VPWR VPWR _17109_/Y sky130_fd_sc_hd__nand2_4
X_18089_ _18089_/A VGND VGND VPWR VPWR _18089_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20120_ _20054_/X _20119_/X _13665_/A _23084_/Q _20117_/X VGND VGND VPWR VPWR _20120_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24565__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20051_ _21154_/B _20048_/X _19731_/X _20048_/X VGND VGND VPWR VPWR _23111_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16635__B1 _24118_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23810_ _23624_/CLK _18626_/X HRESETn VGND VGND VPWR VPWR _23810_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_22_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24790_ _24823_/CLK _14291_/X HRESETn VGND VGND VPWR VPWR _24790_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20953_ _21626_/A _20953_/B _20952_/X VGND VGND VPWR VPWR _20953_/X sky130_fd_sc_hd__and3_4
XFILLER_54_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23741_ _24259_/CLK _20620_/X HRESETn VGND VGND VPWR VPWR _20617_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_96_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20884_ _12062_/X _20882_/X _13326_/A _20883_/X VGND VGND VPWR VPWR _20884_/X sky130_fd_sc_hd__a211o_4
XPHY_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23672_ _23680_/CLK _20371_/Y HRESETn VGND VGND VPWR VPWR _20368_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22623_ _16508_/Y _22435_/X VGND VGND VPWR VPWR _22623_/X sky130_fd_sc_hd__and2_4
XANTENNA__13621__B1 _13330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22554_ _22730_/A _22554_/B VGND VGND VPWR VPWR _22573_/C sky130_fd_sc_hd__nor2_4
XFILLER_42_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21113__D _21275_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21505_ _21374_/A _21505_/B VGND VGND VPWR VPWR _21505_/X sky130_fd_sc_hd__or2_4
XANTENNA__15896__A _24400_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22485_ _20917_/X _22483_/X _20903_/X _22484_/X VGND VGND VPWR VPWR _22486_/B sky130_fd_sc_hd__o22a_4
XFILLER_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21436_ _21300_/A _24258_/Q _13613_/A VGND VGND VPWR VPWR _21436_/X sky130_fd_sc_hd__o21a_4
X_24224_ _24192_/CLK _16384_/X HRESETn VGND VGND VPWR VPWR _16383_/A sky130_fd_sc_hd__dfrtp_4
X_24155_ _24098_/CLK _16571_/X HRESETn VGND VGND VPWR VPWR _24155_/Q sky130_fd_sc_hd__dfrtp_4
X_21367_ _21367_/A _19500_/Y VGND VGND VPWR VPWR _21369_/B sky130_fd_sc_hd__or2_4
X_20318_ _18617_/A _18617_/B VGND VGND VPWR VPWR _20318_/Y sky130_fd_sc_hd__nand2_4
X_23106_ _23109_/CLK _23106_/D VGND VGND VPWR VPWR _20062_/A sky130_fd_sc_hd__dfxtp_4
X_24086_ _24064_/CLK _16867_/X HRESETn VGND VGND VPWR VPWR _24086_/Q sky130_fd_sc_hd__dfrtp_4
X_21298_ _14747_/A _21298_/B VGND VGND VPWR VPWR _21302_/B sky130_fd_sc_hd__or2_4
XFILLER_104_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23037_ _18011_/Y _21491_/A _17224_/Y _23906_/Q VGND VGND VPWR VPWR _23037_/X sky130_fd_sc_hd__a2bb2o_4
X_20249_ _20249_/A _20249_/B VGND VGND VPWR VPWR _20249_/X sky130_fd_sc_hd__and2_4
XFILLER_103_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16626__B1 _24123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24235__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21138__A _21153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14810_ _15003_/A _24147_/Q _15003_/A _24147_/Q VGND VGND VPWR VPWR _14811_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15136__A _15159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19831__A _19831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15790_ _12816_/Y _15787_/X _15511_/X _15787_/X VGND VGND VPWR VPWR _15790_/X sky130_fd_sc_hd__a2bb2o_4
X_24988_ _24953_/CLK _24988_/D HRESETn VGND VGND VPWR VPWR _13353_/A sky130_fd_sc_hd__dfrtp_4
X_14741_ _24711_/Q _14740_/A _14990_/A _14740_/Y VGND VGND VPWR VPWR _14749_/B sky130_fd_sc_hd__o22a_4
X_11953_ _11952_/X VGND VGND VPWR VPWR _11954_/A sky130_fd_sc_hd__buf_2
XFILLER_123_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23939_ _23939_/CLK _23939_/D HRESETn VGND VGND VPWR VPWR _23939_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17460_ _17447_/Y _17460_/B _17459_/Y VGND VGND VPWR VPWR _17460_/X sky130_fd_sc_hd__and3_4
X_14672_ _14657_/X _14671_/Y _24869_/Q _14622_/X VGND VGND VPWR VPWR _14672_/X sky130_fd_sc_hd__a2bb2o_4
X_11884_ _11884_/A _11884_/B VGND VGND VPWR VPWR _11884_/X sky130_fd_sc_hd__and2_4
X_16411_ _24215_/Q VGND VGND VPWR VPWR _16411_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13623_ _11505_/A VGND VGND VPWR VPWR _16043_/A sky130_fd_sc_hd__buf_2
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17391_ _17382_/C _17382_/D VGND VGND VPWR VPWR _17392_/C sky130_fd_sc_hd__nand2_4
XANTENNA__23870__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12495__A _12495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19879__B1 _19835_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25094__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_231_0_HCLK clkbuf_8_231_0_HCLK/A VGND VGND VPWR VPWR _24182_/CLK sky130_fd_sc_hd__clkbuf_1
X_19130_ _19137_/A VGND VGND VPWR VPWR _19130_/X sky130_fd_sc_hd__buf_2
X_16342_ _16341_/Y _16339_/X _16264_/X _16339_/X VGND VGND VPWR VPWR _24240_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13554_ _11676_/Y _11683_/Y VGND VGND VPWR VPWR _13555_/B sky130_fd_sc_hd__or2_4
XFILLER_34_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25023__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12505_ _12505_/A _12505_/B VGND VGND VPWR VPWR _12508_/B sky130_fd_sc_hd__or2_4
X_19061_ _17719_/B VGND VGND VPWR VPWR _19061_/Y sky130_fd_sc_hd__inv_2
X_16273_ _16268_/X _16269_/X _15499_/X _24269_/Q _16270_/X VGND VGND VPWR VPWR _24269_/D
+ sky130_fd_sc_hd__a32o_4
X_13485_ _13468_/Y _13480_/X _13484_/X _21696_/A _13482_/Y VGND VGND VPWR VPWR _24970_/D
+ sky130_fd_sc_hd__a32o_4
X_18012_ _18011_/Y _18008_/X _16671_/X _18008_/X VGND VGND VPWR VPWR _23907_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22416__B _22416_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15224_ _15224_/A _15224_/B VGND VGND VPWR VPWR _15226_/A sky130_fd_sc_hd__nand2_4
X_12436_ _12435_/X VGND VGND VPWR VPWR _25098_/D sky130_fd_sc_hd__inv_2
XFILLER_12_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15155_ _15115_/X _15123_/X _15136_/C VGND VGND VPWR VPWR _15156_/C sky130_fd_sc_hd__o21a_4
X_12367_ _12413_/A VGND VGND VPWR VPWR _12498_/A sky130_fd_sc_hd__buf_2
XFILLER_5_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14106_ _24853_/Q _14106_/B VGND VGND VPWR VPWR _14106_/X sky130_fd_sc_hd__and2_4
XFILLER_5_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16727__A2_N _22395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12298_ _12298_/A VGND VGND VPWR VPWR _12299_/B sky130_fd_sc_hd__inv_2
X_15086_ _15092_/A _15085_/X VGND VGND VPWR VPWR _15093_/B sky130_fd_sc_hd__or2_4
X_19963_ HWDATA[1] VGND VGND VPWR VPWR _19963_/X sky130_fd_sc_hd__buf_2
XFILLER_4_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14037_ _20396_/A _14037_/B VGND VGND VPWR VPWR _14037_/X sky130_fd_sc_hd__or2_4
X_18914_ _18912_/Y _18913_/X _18823_/X _18913_/X VGND VGND VPWR VPWR _18914_/X sky130_fd_sc_hd__a2bb2o_4
X_19894_ _19894_/A VGND VGND VPWR VPWR _21513_/B sky130_fd_sc_hd__inv_2
XFILLER_80_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18845_ _18832_/Y VGND VGND VPWR VPWR _18845_/X sky130_fd_sc_hd__buf_2
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18776_ _18776_/A VGND VGND VPWR VPWR _18776_/X sky130_fd_sc_hd__buf_2
X_15988_ _15986_/Y _15987_/X _15894_/X _15987_/X VGND VGND VPWR VPWR _24366_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22166__A1 _24403_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20887__A _23042_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16284__A1_N _14916_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17727_ _17727_/A VGND VGND VPWR VPWR _17816_/A sky130_fd_sc_hd__buf_2
X_14939_ _24662_/Q VGND VGND VPWR VPWR _14939_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23958__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_41_0_HCLK clkbuf_6_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_83_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17658_ _17657_/Y _15807_/X _17655_/X VGND VGND VPWR VPWR _17658_/X sky130_fd_sc_hd__a21o_4
X_16609_ _16608_/Y _16606_/X _16369_/X _16606_/X VGND VGND VPWR VPWR _16609_/X sky130_fd_sc_hd__a2bb2o_4
X_17589_ _17492_/D _17594_/B VGND VGND VPWR VPWR _17590_/A sky130_fd_sc_hd__or2_4
X_19328_ _19327_/Y VGND VGND VPWR VPWR _19328_/X sky130_fd_sc_hd__buf_2
X_19259_ _16043_/A _23763_/Q _13630_/C _22024_/B VGND VGND VPWR VPWR _19260_/A sky130_fd_sc_hd__and4_4
XANTENNA__15356__B1 _11566_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22270_ _22263_/X _22270_/B VGND VGND VPWR VPWR _22270_/Y sky130_fd_sc_hd__nor2_4
X_21221_ _21385_/A _21221_/B VGND VGND VPWR VPWR _21221_/X sky130_fd_sc_hd__or2_4
XANTENNA__24746__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14125__A _13492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16043__C _16041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21152_ _21340_/A _20112_/Y VGND VGND VPWR VPWR _21152_/X sky130_fd_sc_hd__or2_4
X_20103_ _20110_/A VGND VGND VPWR VPWR _20103_/X sky130_fd_sc_hd__buf_2
XFILLER_8_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21083_ _11960_/A VGND VGND VPWR VPWR _21083_/X sky130_fd_sc_hd__buf_2
XFILLER_99_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20034_ _20034_/A _19644_/X _18031_/C VGND VGND VPWR VPWR _20035_/A sky130_fd_sc_hd__or3_4
XFILLER_119_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24911_ _24904_/CLK _24911_/D HRESETn VGND VGND VPWR VPWR _13818_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_123_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_247_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16623__A3 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24842_ _24962_/CLK _24842_/D HRESETn VGND VGND VPWR VPWR _24842_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14095__B1 _14094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23699__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24773_ _24776_/CLK _14345_/X HRESETn VGND VGND VPWR VPWR _24773_/Q sky130_fd_sc_hd__dfrtp_4
X_21985_ _16202_/A _21984_/X VGND VGND VPWR VPWR _21985_/X sky130_fd_sc_hd__or2_4
XFILLER_2_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21904__B2 _20832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23724_ _24185_/CLK _20544_/X HRESETn VGND VGND VPWR VPWR _20542_/A sky130_fd_sc_hd__dfrtp_4
X_20936_ _21280_/A VGND VGND VPWR VPWR _22011_/A sky130_fd_sc_hd__buf_2
XPHY_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _16473_/Y _21882_/A _24093_/Q _21297_/A VGND VGND VPWR VPWR _20867_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15595__B1 _24528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23655_ _24728_/CLK _23655_/D HRESETn VGND VGND VPWR VPWR _23655_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22606_ _22178_/A VGND VGND VPWR VPWR _22606_/X sky130_fd_sc_hd__buf_2
X_20798_ _22870_/B VGND VGND VPWR VPWR _22148_/A sky130_fd_sc_hd__buf_2
XPHY_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23586_ _23586_/CLK _18725_/X VGND VGND VPWR VPWR _23586_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22537_ _21544_/A VGND VGND VPWR VPWR _22537_/X sky130_fd_sc_hd__buf_2
XFILLER_22_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_61_0_HCLK clkbuf_7_30_0_HCLK/X VGND VGND VPWR VPWR _23972_/CLK sky130_fd_sc_hd__clkbuf_1
X_13270_ _13238_/A _13270_/B _13270_/C VGND VGND VPWR VPWR _13271_/C sky130_fd_sc_hd__and3_4
X_22468_ _22468_/A VGND VGND VPWR VPWR _22468_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11908__B1 _11904_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12221_ _12207_/B VGND VGND VPWR VPWR _12222_/B sky130_fd_sc_hd__inv_2
XANTENNA__18297__C1 _18228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24487__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24207_ _23830_/CLK _16431_/X HRESETn VGND VGND VPWR VPWR _24207_/Q sky130_fd_sc_hd__dfrtp_4
X_21419_ _16467_/A _22155_/A VGND VGND VPWR VPWR _21422_/B sky130_fd_sc_hd__or2_4
X_22399_ _22399_/A _22312_/B VGND VGND VPWR VPWR _22399_/Y sky130_fd_sc_hd__nor2_4
X_25187_ _23353_/CLK _11715_/X HRESETn VGND VGND VPWR VPWR _11698_/D sky130_fd_sc_hd__dfrtp_4
X_12152_ _12152_/A VGND VGND VPWR VPWR _12152_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24416__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24138_ _24138_/CLK _16599_/X HRESETn VGND VGND VPWR VPWR _24138_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_2_2_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12083_ _12083_/A VGND VGND VPWR VPWR _12083_/X sky130_fd_sc_hd__buf_2
X_16960_ _16133_/Y _24058_/Q _16133_/Y _24058_/Q VGND VGND VPWR VPWR _16960_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_123_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24069_ _24623_/CLK _24069_/D HRESETn VGND VGND VPWR VPWR _16758_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_2_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12333__B1 _12448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15911_ _11535_/X _15641_/X _15735_/X _20737_/A _15910_/X VGND VGND VPWR VPWR _24394_/D
+ sky130_fd_sc_hd__a32o_4
X_16891_ _16800_/Y _16885_/X _16858_/X _16888_/B VGND VGND VPWR VPWR _16891_/X sky130_fd_sc_hd__a211o_4
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18630_ _18607_/A _18620_/Y _23644_/Q _20705_/B _18624_/A VGND VGND VPWR VPWR _23806_/D
+ sky130_fd_sc_hd__a32o_4
X_15842_ _15847_/A VGND VGND VPWR VPWR _15842_/X sky130_fd_sc_hd__buf_2
XFILLER_65_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16614__A3 _15706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18561_ pwm_S7 VGND VGND VPWR VPWR _18561_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15773_ _15767_/X VGND VGND VPWR VPWR _15773_/X sky130_fd_sc_hd__buf_2
X_12985_ _12815_/Y _12984_/X _12896_/X VGND VGND VPWR VPWR _12985_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_79_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17512_ _17505_/B _17511_/X VGND VGND VPWR VPWR _17512_/X sky130_fd_sc_hd__or2_4
XFILLER_79_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14724_ _24690_/Q VGND VGND VPWR VPWR _14872_/B sky130_fd_sc_hd__inv_2
Xclkbuf_5_28_0_HCLK clkbuf_4_14_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_11936_ _25156_/Q VGND VGND VPWR VPWR _11936_/Y sky130_fd_sc_hd__inv_2
X_18492_ _18504_/A _18492_/B _18492_/C VGND VGND VPWR VPWR _18492_/X sky130_fd_sc_hd__and3_4
XFILLER_75_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18772__B1 _18700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25204__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17443_ _17434_/X _17443_/B _17428_/C VGND VGND VPWR VPWR _17443_/X sky130_fd_sc_hd__and3_4
X_14655_ _14655_/A VGND VGND VPWR VPWR _14655_/X sky130_fd_sc_hd__buf_2
XANTENNA__15586__B1 _24533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11867_ _11868_/A _11866_/X VGND VGND VPWR VPWR _11867_/X sky130_fd_sc_hd__and2_4
XFILLER_60_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13606_ _11683_/A _13594_/X _13576_/X _11683_/Y VGND VGND VPWR VPWR _24947_/D sky130_fd_sc_hd__o22a_4
X_17374_ _17373_/X VGND VGND VPWR VPWR _17375_/B sky130_fd_sc_hd__inv_2
X_14586_ _18873_/B VGND VGND VPWR VPWR _19946_/A sky130_fd_sc_hd__inv_2
X_11798_ _11772_/B _11796_/Y _11797_/Y VGND VGND VPWR VPWR _11798_/X sky130_fd_sc_hd__o21a_4
X_19113_ _23449_/Q VGND VGND VPWR VPWR _19113_/Y sky130_fd_sc_hd__inv_2
X_16325_ _16325_/A VGND VGND VPWR VPWR _16325_/Y sky130_fd_sc_hd__inv_2
X_13537_ _20656_/A _20653_/B _13537_/C VGND VGND VPWR VPWR _13537_/X sky130_fd_sc_hd__or3_4
XANTENNA__15338__B1 _11545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22146__B _22146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19044_ _23475_/Q VGND VGND VPWR VPWR _19044_/Y sky130_fd_sc_hd__inv_2
X_16256_ _16256_/A VGND VGND VPWR VPWR _16262_/A sky130_fd_sc_hd__buf_2
XANTENNA__20882__B2 _11527_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13468_ _13468_/A _13468_/B VGND VGND VPWR VPWR _13468_/Y sky130_fd_sc_hd__nand2_4
X_15207_ _15192_/A _15207_/B _15207_/C VGND VGND VPWR VPWR _15207_/X sky130_fd_sc_hd__and3_4
X_12419_ _12419_/A VGND VGND VPWR VPWR _12419_/Y sky130_fd_sc_hd__inv_2
X_16187_ _16186_/Y _16184_/X _16093_/X _16184_/X VGND VGND VPWR VPWR _24302_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13399_ SSn_S2 _13397_/Y _13398_/X _13397_/Y VGND VGND VPWR VPWR _24974_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24157__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15138_ _15138_/A _15138_/B _14898_/Y _15154_/B VGND VGND VPWR VPWR _15139_/A sky130_fd_sc_hd__or4_4
XFILLER_126_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14313__A1 _23077_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15069_ _15068_/X VGND VGND VPWR VPWR _24692_/D sky130_fd_sc_hd__inv_2
X_19946_ _19946_/A _19946_/B _19946_/C _19100_/B VGND VGND VPWR VPWR _19946_/X sky130_fd_sc_hd__or4_4
XANTENNA__15510__B1 _13658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19877_ _21392_/B _19876_/X _19832_/X _19876_/X VGND VGND VPWR VPWR _19877_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19252__B2 _19251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18828_ _18711_/X VGND VGND VPWR VPWR _18828_/X sky130_fd_sc_hd__buf_2
XFILLER_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15813__A1 _16222_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22139__B2 _20927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13008__B _13008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23792__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18759_ _14587_/A _18759_/B _13461_/X VGND VGND VPWR VPWR _18760_/A sky130_fd_sc_hd__or3_4
XFILLER_82_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15504__A _15460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21770_ _21762_/X _18837_/Y VGND VGND VPWR VPWR _21771_/C sky130_fd_sc_hd__or2_4
XANTENNA__23721__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20721_ scl_oen_o_S5 _20720_/Y VGND VGND VPWR VPWR _20721_/X sky130_fd_sc_hd__and2_4
XFILLER_19_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20652_ _20647_/X _20650_/X _24179_/Q _20651_/X VGND VGND VPWR VPWR _23748_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24998__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23440_ _23440_/CLK _19140_/X VGND VGND VPWR VPWR _23440_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13052__B2 _11708_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21241__A _21394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24927__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23371_ _23374_/CLK _19337_/X VGND VGND VPWR VPWR _23371_/Q sky130_fd_sc_hd__dfxtp_4
X_20583_ _20555_/A VGND VGND VPWR VPWR _20583_/X sky130_fd_sc_hd__buf_2
XFILLER_109_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_48_0_HCLK clkbuf_7_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_48_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_25110_ _25115_/CLK _25110_/D HRESETn VGND VGND VPWR VPWR _12097_/A sky130_fd_sc_hd__dfrtp_4
X_22322_ _22322_/A VGND VGND VPWR VPWR _22322_/X sky130_fd_sc_hd__buf_2
XANTENNA__20873__B2 _15426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_19_0_HCLK_A clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22253_ _20748_/X _22248_/Y _21029_/X _22252_/X VGND VGND VPWR VPWR _22254_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24580__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25041_ _25067_/CLK _25041_/D HRESETn VGND VGND VPWR VPWR _25041_/Q sky130_fd_sc_hd__dfrtp_4
X_21204_ _21374_/A _19461_/Y VGND VGND VPWR VPWR _21207_/B sky130_fd_sc_hd__or2_4
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22184_ _12346_/A _22153_/B VGND VGND VPWR VPWR _22184_/X sky130_fd_sc_hd__or2_4
X_21135_ _21130_/X _21132_/X _21134_/X VGND VGND VPWR VPWR _21135_/X sky130_fd_sc_hd__and3_4
XFILLER_8_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21075__A2_N _12062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16070__A _24345_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22378__B2 _22121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21066_ _21066_/A _21066_/B VGND VGND VPWR VPWR _21066_/X sky130_fd_sc_hd__and2_4
XFILLER_119_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22917__A3 _22839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20017_ _23124_/Q VGND VGND VPWR VPWR _21917_/B sky130_fd_sc_hd__inv_2
XANTENNA__19381__A _11625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17254__B1 _11606_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15804__A1 _15799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15804__B2 _15746_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24825_ _24851_/CLK _24825_/D HRESETn VGND VGND VPWR VPWR _24825_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12618__B2 _12617_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15414__A _15414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12770_ _12650_/A _12770_/B VGND VGND VPWR VPWR _12770_/X sky130_fd_sc_hd__or2_4
XPHY_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24756_ _24757_/CLK _24756_/D HRESETn VGND VGND VPWR VPWR _14420_/A sky130_fd_sc_hd__dfrtp_4
X_21968_ _20940_/X _21923_/X _21938_/X _20918_/X _21967_/Y VGND VGND VPWR VPWR _21968_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22550__A1 _14838_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22550__B2 _22549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _24618_/Q VGND VGND VPWR VPWR _14013_/A sky130_fd_sc_hd__inv_2
XFILLER_37_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23707_ _23706_/CLK _23707_/D HRESETn VGND VGND VPWR VPWR _13508_/D sky130_fd_sc_hd__dfrtp_4
X_20919_ _20919_/A _20866_/X VGND VGND VPWR VPWR _20919_/X sky130_fd_sc_hd__and2_4
XPHY_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24687_ _24674_/CLK _15082_/X HRESETn VGND VGND VPWR VPWR _24687_/Q sky130_fd_sc_hd__dfrtp_4
X_21899_ _22006_/B _21897_/X _21881_/A _21898_/X VGND VGND VPWR VPWR _21899_/X sky130_fd_sc_hd__o22a_4
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _24745_/Q VGND VGND VPWR VPWR _14440_/X sky130_fd_sc_hd__buf_2
XFILLER_120_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _13557_/A _23914_/Q _13564_/A _11665_/A VGND VGND VPWR VPWR _11652_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23638_ _24811_/CLK _20317_/Y HRESETn VGND VGND VPWR VPWR _18616_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14240__B1 _14209_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21151__A _17629_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24668__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14371_ _14390_/D VGND VGND VPWR VPWR _14371_/X sky130_fd_sc_hd__buf_2
XPHY_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11583_ _11583_/A VGND VGND VPWR VPWR _11583_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16759__A1_N _24405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23569_ _23568_/CLK _23569_/D VGND VGND VPWR VPWR _23569_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16110_ _22014_/A _16105_/X _15890_/X _16105_/X VGND VGND VPWR VPWR _16110_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13322_ _23041_/A VGND VGND VPWR VPWR _20891_/A sky130_fd_sc_hd__inv_2
XFILLER_35_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17090_ _17101_/A _17077_/X _17090_/C VGND VGND VPWR VPWR _17090_/X sky130_fd_sc_hd__and3_4
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16041_ _21273_/A VGND VGND VPWR VPWR _16041_/X sky130_fd_sc_hd__buf_2
X_13253_ _13221_/A _13251_/X _13253_/C VGND VGND VPWR VPWR _13254_/C sky130_fd_sc_hd__and3_4
XFILLER_129_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12204_ _12170_/B _12193_/B _12203_/X _12200_/B VGND VGND VPWR VPWR _12204_/X sky130_fd_sc_hd__a211o_4
XFILLER_108_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24250__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_5_0_HCLK clkbuf_6_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13184_ _13102_/X _13182_/X _13183_/X VGND VGND VPWR VPWR _13184_/X sky130_fd_sc_hd__and3_4
X_19800_ _19801_/A VGND VGND VPWR VPWR _19800_/X sky130_fd_sc_hd__buf_2
X_12135_ _12207_/A _24568_/Q _12207_/A _24568_/Q VGND VGND VPWR VPWR _12140_/B sky130_fd_sc_hd__a2bb2o_4
X_17992_ _11680_/Y _17987_/X _16455_/X _17987_/X VGND VGND VPWR VPWR _23918_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12306__B1 _12305_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16943_ _24064_/Q _16942_/Y VGND VGND VPWR VPWR _16943_/X sky130_fd_sc_hd__or2_4
X_19731_ _11855_/A VGND VGND VPWR VPWR _19731_/X sky130_fd_sc_hd__buf_2
X_12066_ _16559_/A VGND VGND VPWR VPWR _16302_/A sky130_fd_sc_hd__buf_2
XFILLER_104_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14212__B _14199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13109__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16874_ _16769_/Y _16874_/B VGND VGND VPWR VPWR _16874_/Y sky130_fd_sc_hd__nand2_4
X_19662_ _19661_/Y _19659_/X _19617_/X _19659_/X VGND VGND VPWR VPWR _23256_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15825_ _15824_/X VGND VGND VPWR VPWR _15826_/A sky130_fd_sc_hd__buf_2
X_18613_ _20301_/A _20298_/A VGND VGND VPWR VPWR _18614_/B sky130_fd_sc_hd__or2_4
XFILLER_93_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19593_ _21013_/B _19588_/X _19506_/X _19575_/Y VGND VGND VPWR VPWR _19593_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11852__A _11830_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15756_ HWDATA[27] VGND VGND VPWR VPWR _15756_/X sky130_fd_sc_hd__buf_2
X_18544_ _18540_/A _18535_/B _18544_/C VGND VGND VPWR VPWR _23819_/D sky130_fd_sc_hd__and3_4
X_12968_ _12992_/A _12966_/X _12967_/X VGND VGND VPWR VPWR _25018_/D sky130_fd_sc_hd__and3_4
XFILLER_64_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14707_ _14876_/D VGND VGND VPWR VPWR _15033_/A sky130_fd_sc_hd__buf_2
X_11919_ _11919_/A VGND VGND VPWR VPWR _11919_/X sky130_fd_sc_hd__buf_2
X_18475_ _18475_/A VGND VGND VPWR VPWR _18475_/X sky130_fd_sc_hd__buf_2
X_15687_ _15684_/X _15672_/X _16087_/A _24482_/Q _15685_/X VGND VGND VPWR VPWR _15687_/X
+ sky130_fd_sc_hd__a32o_4
X_12899_ _12963_/A _12885_/X _12899_/C _12779_/Y VGND VGND VPWR VPWR _12899_/X sky130_fd_sc_hd__or4_4
XFILLER_127_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17426_ _17317_/D _17411_/B VGND VGND VPWR VPWR _17426_/Y sky130_fd_sc_hd__nand2_4
X_14638_ _24729_/Q _14615_/A _14608_/Y _14615_/Y VGND VGND VPWR VPWR _14638_/X sky130_fd_sc_hd__o22a_4
XFILLER_14_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17357_ _17356_/X VGND VGND VPWR VPWR _24004_/D sky130_fd_sc_hd__inv_2
X_14569_ _14569_/A VGND VGND VPWR VPWR _17702_/A sky130_fd_sc_hd__buf_2
XFILLER_119_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16308_ _16308_/A VGND VGND VPWR VPWR _16308_/X sky130_fd_sc_hd__buf_2
XANTENNA__24338__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17288_ _24000_/Q VGND VGND VPWR VPWR _17288_/Y sky130_fd_sc_hd__inv_2
X_19027_ _19027_/A VGND VGND VPWR VPWR _21209_/B sky130_fd_sc_hd__inv_2
X_16239_ _16228_/X _16234_/X _15468_/X _24285_/Q _16237_/X VGND VGND VPWR VPWR _24285_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14298__B1 _14221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19929_ _19929_/A VGND VGND VPWR VPWR _21943_/B sky130_fd_sc_hd__inv_2
XFILLER_130_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23021__A2 _22859_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23973__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25197__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23902__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22940_ _11524_/Y _22536_/X _15927_/Y _22537_/X VGND VGND VPWR VPWR _22940_/X sky130_fd_sc_hd__o22a_4
XFILLER_112_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25126__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15798__B1 _15279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22871_ _21864_/X _22869_/X _22530_/X _22870_/X VGND VGND VPWR VPWR _22871_/X sky130_fd_sc_hd__o22a_4
X_24610_ _24185_/CLK _15338_/X HRESETn VGND VGND VPWR VPWR _24610_/Q sky130_fd_sc_hd__dfrtp_4
X_21822_ _20978_/A _19693_/Y VGND VGND VPWR VPWR _21825_/B sky130_fd_sc_hd__or2_4
XFILLER_37_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22532__B2 _22531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_11_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_24541_ _23179_/CLK _15538_/X HRESETn VGND VGND VPWR VPWR _24541_/Q sky130_fd_sc_hd__dfrtp_4
X_21753_ _24749_/Q _19273_/Y _21750_/X _21752_/X VGND VGND VPWR VPWR _21753_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20704_ _13950_/A _20703_/X _13923_/B VGND VGND VPWR VPWR _20704_/X sky130_fd_sc_hd__o21a_4
XFILLER_58_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24472_ _24307_/CLK _15703_/X HRESETn VGND VGND VPWR VPWR _24472_/Q sky130_fd_sc_hd__dfrtp_4
X_21684_ _21009_/A VGND VGND VPWR VPWR _22064_/A sky130_fd_sc_hd__buf_2
XANTENNA__14222__B1 _14221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22067__A _21396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24761__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23423_ _23425_/CLK _23423_/D VGND VGND VPWR VPWR _17949_/B sky130_fd_sc_hd__dfxtp_4
X_20635_ _20635_/A _20635_/B _20635_/C _20653_/A VGND VGND VPWR VPWR _20635_/X sky130_fd_sc_hd__or4_4
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24079__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20566_ _23730_/Q VGND VGND VPWR VPWR _20566_/Y sky130_fd_sc_hd__inv_2
X_23354_ _23336_/CLK _19384_/X VGND VGND VPWR VPWR _13216_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_20_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24008__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22305_ _20748_/X _22302_/Y _21029_/X _22304_/X VGND VGND VPWR VPWR _22305_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22048__B1 _24932_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20497_ _20484_/X _20496_/Y _15361_/A _20488_/X VGND VGND VPWR VPWR _23712_/D sky130_fd_sc_hd__a2bb2o_4
X_23285_ _23282_/CLK _23285_/D VGND VGND VPWR VPWR _23285_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22599__A1 _22369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25024_ _25021_/CLK _25024_/D HRESETn VGND VGND VPWR VPWR _22651_/A sky130_fd_sc_hd__dfrtp_4
X_22236_ _22201_/X _22205_/X _22209_/X _22222_/Y _22235_/Y VGND VGND VPWR VPWR HRDATA[9]
+ sky130_fd_sc_hd__a2111o_4
Xclkbuf_8_135_0_HCLK clkbuf_7_67_0_HCLK/X VGND VGND VPWR VPWR _23419_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_106_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_198_0_HCLK clkbuf_7_99_0_HCLK/X VGND VGND VPWR VPWR _23734_/CLK sky130_fd_sc_hd__clkbuf_1
X_22167_ _22167_/A _22164_/X _22167_/C VGND VGND VPWR VPWR _22168_/C sky130_fd_sc_hd__and3_4
XANTENNA__15409__A _21113_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14289__B1 _14228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21118_ _12054_/A _20872_/X _18127_/Y _11960_/A VGND VGND VPWR VPWR _21118_/X sky130_fd_sc_hd__o22a_4
X_22098_ _17636_/A _22090_/X _22097_/X VGND VGND VPWR VPWR _22114_/C sky130_fd_sc_hd__and3_4
XANTENNA__22530__A _22610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21023__A1 _13624_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13940_ _13998_/B _13926_/B _24884_/Q VGND VGND VPWR VPWR _13941_/B sky130_fd_sc_hd__or3_4
X_21049_ _21049_/A VGND VGND VPWR VPWR _21049_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17624__A _17460_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23643__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21574__A2 _21553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22771__A1 _17481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16053__A1_N _16050_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21146__A _21336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13871_ _13808_/X _13810_/X _13811_/A _13806_/X VGND VGND VPWR VPWR _13871_/X sky130_fd_sc_hd__or4_4
XANTENNA__15789__B1 _15788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15610_ _12592_/Y _15607_/X _11573_/X _15607_/X VGND VGND VPWR VPWR _24519_/D sky130_fd_sc_hd__a2bb2o_4
X_12822_ _12783_/X _12822_/B _12808_/X _12821_/X VGND VGND VPWR VPWR _12822_/X sky130_fd_sc_hd__or4_4
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24808_ _24788_/CLK _14246_/X HRESETn VGND VGND VPWR VPWR _14009_/A sky130_fd_sc_hd__dfstp_4
X_16590_ _16566_/A VGND VGND VPWR VPWR _16590_/X sky130_fd_sc_hd__buf_2
XANTENNA__20129__A3 _11643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15541_ _19442_/A VGND VGND VPWR VPWR _15541_/X sky130_fd_sc_hd__buf_2
XANTENNA__24849__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12753_ _12749_/A _12741_/B _12753_/C VGND VGND VPWR VPWR _25044_/D sky130_fd_sc_hd__and3_4
XPHY_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24739_ _24740_/CLK _24739_/D HRESETn VGND VGND VPWR VPWR _24739_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11703_/X VGND VGND VPWR VPWR _11704_/Y sky130_fd_sc_hd__inv_2
X_18260_ _18559_/B _18260_/B _18259_/X VGND VGND VPWR VPWR _18260_/X sky130_fd_sc_hd__or3_4
XFILLER_37_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ _15472_/A VGND VGND VPWR VPWR _15472_/X sky130_fd_sc_hd__buf_2
XFILLER_91_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12727_/A _12655_/X _12679_/C VGND VGND VPWR VPWR _12685_/C sky130_fd_sc_hd__o21a_4
XPHY_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17210_/Y _17206_/X _16211_/X _17206_/X VGND VGND VPWR VPWR _17211_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14374_/X _14422_/Y _14371_/X _14415_/X _13447_/A VGND VGND VPWR VPWR _24755_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ _11635_/A VGND VGND VPWR VPWR _15801_/A sky130_fd_sc_hd__buf_2
X_18191_ _18172_/X _18191_/B _18191_/C _18190_/X VGND VGND VPWR VPWR _18192_/B sky130_fd_sc_hd__or4_4
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17142_ _16966_/Y _17141_/X _17074_/A _17137_/B VGND VGND VPWR VPWR _17143_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24431__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14354_ scl_oen_o_S4 _14348_/X _14349_/Y _14353_/Y VGND VGND VPWR VPWR _14355_/B
+ sky130_fd_sc_hd__o22a_4
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11566_ HWDATA[19] VGND VGND VPWR VPWR _11566_/X sky130_fd_sc_hd__buf_2
XFILLER_7_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13305_ _13204_/A _13305_/B VGND VGND VPWR VPWR _13307_/B sky130_fd_sc_hd__or2_4
Xclkbuf_7_31_0_HCLK clkbuf_7_30_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17073_ _17045_/X _17054_/B _17023_/Y VGND VGND VPWR VPWR _17073_/X sky130_fd_sc_hd__o21a_4
XFILLER_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14285_ _14284_/Y _14280_/X _14218_/X _14273_/A VGND VGND VPWR VPWR _24792_/D sky130_fd_sc_hd__a2bb2o_4
X_11497_ _24618_/Q VGND VGND VPWR VPWR _11938_/A sky130_fd_sc_hd__buf_2
XFILLER_13_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22424__B _11964_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_94_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_94_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_16024_ _16023_/X VGND VGND VPWR VPWR _16024_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13236_ _13300_/A _23601_/Q VGND VGND VPWR VPWR _13238_/B sky130_fd_sc_hd__or2_4
XFILLER_40_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20065__A2 _15410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15319__A _15531_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11847__A _19610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13167_ _13203_/A _13167_/B _13166_/X VGND VGND VPWR VPWR _13172_/B sky130_fd_sc_hd__and3_4
XFILLER_135_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16636__A1_N _14729_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14819__A2 _14818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12118_ _12116_/A _12117_/A _12174_/A _12117_/Y VGND VGND VPWR VPWR _12118_/X sky130_fd_sc_hd__o22a_4
X_13098_ _13016_/A VGND VGND VPWR VPWR _13316_/A sky130_fd_sc_hd__buf_2
X_17975_ _17974_/X VGND VGND VPWR VPWR _17975_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17218__B1 _16556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_HCLK clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19714_ _19714_/A VGND VGND VPWR VPWR _19714_/X sky130_fd_sc_hd__buf_2
X_12049_ _12049_/A _12048_/X VGND VGND VPWR VPWR _12051_/A sky130_fd_sc_hd__or2_4
X_16926_ _16935_/A _16938_/B VGND VGND VPWR VPWR _16936_/B sky130_fd_sc_hd__or2_4
XFILLER_78_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21056__A _21034_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19645_ _18020_/X _18039_/X _20034_/A _19644_/X VGND VGND VPWR VPWR _19646_/A sky130_fd_sc_hd__or4_4
XFILLER_4_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16857_ _16867_/A _16855_/X _16856_/X VGND VGND VPWR VPWR _24088_/D sky130_fd_sc_hd__and3_4
XFILLER_65_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15808_ _16222_/C _15806_/Y _15807_/X VGND VGND VPWR VPWR _15808_/X sky130_fd_sc_hd__o21a_4
X_16788_ _24396_/Q _16921_/C _24400_/Q _16923_/A VGND VGND VPWR VPWR _16791_/B sky130_fd_sc_hd__a2bb2o_4
X_19576_ _19575_/Y VGND VGND VPWR VPWR _19576_/X sky130_fd_sc_hd__buf_2
XANTENNA__21317__A2 _15653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15739_ _15411_/X _15617_/X _15735_/X _24462_/Q _15738_/X VGND VGND VPWR VPWR _24462_/D
+ sky130_fd_sc_hd__a32o_4
X_18527_ _18529_/B VGND VGND VPWR VPWR _18527_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24519__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18458_ _18458_/A VGND VGND VPWR VPWR _18458_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17409_ _17321_/Y _17409_/B VGND VGND VPWR VPWR _17429_/A sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_3_5_0_HCLK_A clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18389_ _16416_/Y _18479_/A _16416_/Y _18388_/A VGND VGND VPWR VPWR _18389_/X sky130_fd_sc_hd__a2bb2o_4
X_20420_ _15405_/Y _20416_/X _21020_/A _20419_/X VGND VGND VPWR VPWR _20420_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20828__A1 _24462_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24172__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20828__B2 _20827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22615__A _14737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24101__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20351_ _14057_/Y _20344_/X _20401_/A _20350_/X VGND VGND VPWR VPWR _20352_/A sky130_fd_sc_hd__a211o_4
XFILLER_134_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23070_ _23992_/CLK _20151_/X VGND VGND VPWR VPWR _23070_/Q sky130_fd_sc_hd__dfxtp_4
X_20282_ _23631_/Q _20279_/A VGND VGND VPWR VPWR _20282_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__20135__A _20134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22021_ _22011_/X _22013_/X _22497_/B _22020_/X VGND VGND VPWR VPWR _22022_/A sky130_fd_sc_hd__o22a_4
XFILLER_88_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20056__A2 _15410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_208_0_HCLK clkbuf_7_104_0_HCLK/X VGND VGND VPWR VPWR _24222_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21253__B2 _21720_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22350__A _22616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17209__B1 _16546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23972_ _23972_/CLK _17514_/Y HRESETn VGND VGND VPWR VPWR _22979_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_111_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24802__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22923_ _22982_/A _22920_/X _22921_/X _22923_/D VGND VGND VPWR VPWR _22923_/X sky130_fd_sc_hd__or4_4
XFILLER_21_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24865__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22854_ _22854_/A _22418_/X VGND VGND VPWR VPWR _22854_/X sky130_fd_sc_hd__and2_4
XFILLER_72_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15786__A3 _16100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18709__B1 _18685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16983__A2 _24046_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21805_ _21805_/A _20064_/X VGND VGND VPWR VPWR _21805_/X sky130_fd_sc_hd__and2_4
XANTENNA__24942__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22785_ _22971_/A _22782_/X _22784_/X VGND VGND VPWR VPWR _22785_/X sky130_fd_sc_hd__and3_4
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19382__B1 _19381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24524_ _25005_/CLK _24524_/D HRESETn VGND VGND VPWR VPWR _12619_/A sky130_fd_sc_hd__dfrtp_4
X_21736_ _14052_/Y _21083_/X _20393_/A _21425_/B VGND VGND VPWR VPWR _21737_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24455_ _24478_/CLK _24455_/D HRESETn VGND VGND VPWR VPWR _24455_/Q sky130_fd_sc_hd__dfrtp_4
X_21667_ _21008_/A VGND VGND VPWR VPWR _21667_/X sky130_fd_sc_hd__buf_2
XANTENNA__22808__A2 _21553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23406_ _23246_/CLK _23406_/D VGND VGND VPWR VPWR _23406_/Q sky130_fd_sc_hd__dfxtp_4
X_20618_ _20617_/A _13535_/X VGND VGND VPWR VPWR _20618_/X sky130_fd_sc_hd__or2_4
X_24386_ _24385_/CLK _15937_/X HRESETn VGND VGND VPWR VPWR _22838_/A sky130_fd_sc_hd__dfrtp_4
X_21598_ _21064_/Y _21594_/X _21596_/X _20800_/A _21597_/X VGND VGND VPWR VPWR _21598_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19685__B2 _19680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17696__B1 _16678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_18_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_18_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_23337_ _23336_/CLK _23337_/D VGND VGND VPWR VPWR _13251_/B sky130_fd_sc_hd__dfxtp_4
X_20549_ _20413_/A _23726_/Q _13515_/X _23026_/A _20465_/X VGND VGND VPWR VPWR _23726_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_4_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21492__B2 _15642_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16523__A _16499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14070_ _13794_/A _15251_/A _13800_/A VGND VGND VPWR VPWR _14070_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_10_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19437__B2 _19417_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23895__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23268_ _23242_/CLK _19630_/X VGND VGND VPWR VPWR _23268_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_134_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13021_ _13299_/A VGND VGND VPWR VPWR _13047_/A sky130_fd_sc_hd__buf_2
X_25007_ _25012_/CLK _13004_/X HRESETn VGND VGND VPWR VPWR _25007_/Q sky130_fd_sc_hd__dfrtp_4
X_22219_ _22219_/A VGND VGND VPWR VPWR _22354_/A sky130_fd_sc_hd__buf_2
XFILLER_106_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23824__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23199_ _24005_/CLK _19811_/X VGND VGND VPWR VPWR _23199_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25048__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16120__B1 _15282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22260__A _21434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14972_ _14965_/X _14972_/B _14972_/C _14971_/X VGND VGND VPWR VPWR _14972_/X sky130_fd_sc_hd__or4_4
X_17760_ _14577_/X VGND VGND VPWR VPWR _17903_/A sky130_fd_sc_hd__buf_2
XFILLER_94_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21547__A2 _11986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18948__B1 _18880_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13923_ scl_oen_o_S4 _13923_/B _13923_/C VGND VGND VPWR VPWR _13934_/B sky130_fd_sc_hd__and3_4
X_16711_ _24389_/Q _16710_/A _15927_/Y _16710_/Y VGND VGND VPWR VPWR _16716_/B sky130_fd_sc_hd__o22a_4
X_17691_ _17694_/A _23446_/Q VGND VGND VPWR VPWR _17692_/C sky130_fd_sc_hd__or2_4
XANTENNA__12498__A _12498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16642_ _16628_/A VGND VGND VPWR VPWR _16643_/A sky130_fd_sc_hd__buf_2
X_19430_ _19429_/Y _19425_/X _19360_/X _19425_/X VGND VGND VPWR VPWR _23338_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13854_ _13822_/B _13848_/X _14361_/B VGND VGND VPWR VPWR _13854_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12805_ _22133_/A VGND VGND VPWR VPWR _12805_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24683__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16573_ _16234_/A VGND VGND VPWR VPWR _16573_/X sky130_fd_sc_hd__buf_2
X_19361_ _19359_/Y _19355_/X _19360_/X _19355_/X VGND VGND VPWR VPWR _23362_/D sky130_fd_sc_hd__a2bb2o_4
X_13785_ _13783_/Y _13785_/B _13769_/D _13766_/D VGND VGND VPWR VPWR _13786_/A sky130_fd_sc_hd__or4_4
XFILLER_43_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15524_ _12114_/Y _15518_/X _15286_/X _15518_/X VGND VGND VPWR VPWR _15524_/X sky130_fd_sc_hd__a2bb2o_4
X_18312_ _18312_/A _18312_/B VGND VGND VPWR VPWR _18312_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12996__B1 _12922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22419__B _11964_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24612__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12736_ _12629_/X _12584_/Y _12651_/C _12735_/X VGND VGND VPWR VPWR _12737_/B sky130_fd_sc_hd__or4_4
X_19292_ _21632_/B _19289_/X _11848_/X _19289_/X VGND VGND VPWR VPWR _23387_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16187__B1 _16093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21323__B _21323_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18243_ _18243_/A VGND VGND VPWR VPWR _18248_/B sky130_fd_sc_hd__inv_2
X_15455_ _11950_/X _16038_/B _14195_/C _11514_/A VGND VGND VPWR VPWR _15455_/X sky130_fd_sc_hd__or4_4
XANTENNA__22138__C _22138_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12667_ _12657_/A _12664_/X _12658_/Y _12666_/X VGND VGND VPWR VPWR _12668_/A sky130_fd_sc_hd__a211o_4
XANTENNA__15934__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14218__A _14218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18913__A _18899_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ _14402_/B _14399_/X _14405_/Y _14403_/X _24762_/Q VGND VGND VPWR VPWR _14406_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_15_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11618_ _25195_/Q VGND VGND VPWR VPWR _11618_/Y sky130_fd_sc_hd__inv_2
X_18174_ _16066_/Y _18256_/A _16066_/Y _18256_/A VGND VGND VPWR VPWR _18177_/B sky130_fd_sc_hd__a2bb2o_4
X_15386_ _16369_/A VGND VGND VPWR VPWR _15386_/X sky130_fd_sc_hd__buf_2
X_12598_ _25049_/Q VGND VGND VPWR VPWR _12728_/A sky130_fd_sc_hd__inv_2
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22435__A _20832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17125_ _17043_/B _17124_/X VGND VGND VPWR VPWR _17126_/A sky130_fd_sc_hd__or2_4
XFILLER_89_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14337_ _14335_/X _14336_/X _24789_/Q _14331_/X VGND VGND VPWR VPWR _14337_/X sky130_fd_sc_hd__o22a_4
X_11549_ _11547_/Y _11542_/X _11548_/X _11542_/X VGND VGND VPWR VPWR _11549_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16433__A _16401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22154__B _22154_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17056_ _17086_/A VGND VGND VPWR VPWR _17056_/Y sky130_fd_sc_hd__inv_2
X_14268_ _14273_/A VGND VGND VPWR VPWR _14268_/X sky130_fd_sc_hd__buf_2
XFILLER_100_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16007_ _16005_/X _16006_/X VGND VGND VPWR VPWR _16221_/C sky130_fd_sc_hd__nor2_4
XFILLER_83_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13219_ _13219_/A _19429_/A VGND VGND VPWR VPWR _13219_/X sky130_fd_sc_hd__or2_4
XANTENNA__22432__B1 _21642_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21993__B _22524_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14199_ _13934_/A _14199_/B VGND VGND VPWR VPWR _14201_/A sky130_fd_sc_hd__nor2_4
XFILLER_97_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_181_0_HCLK clkbuf_7_90_0_HCLK/X VGND VGND VPWR VPWR _24459_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22170__A _21020_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_38_0_HCLK clkbuf_8_39_0_HCLK/A VGND VGND VPWR VPWR _23471_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_135_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17958_ _17783_/A _17958_/B _17957_/X VGND VGND VPWR VPWR _17962_/B sky130_fd_sc_hd__and3_4
XANTENNA__18939__B1 _18938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16909_ _16825_/Y _16885_/B _16858_/X _16907_/B VGND VGND VPWR VPWR _16910_/A sky130_fd_sc_hd__a211o_4
X_17889_ _17889_/A _17889_/B _17888_/X VGND VGND VPWR VPWR _17889_/X sky130_fd_sc_hd__and3_4
XFILLER_81_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19628_ _23268_/Q VGND VGND VPWR VPWR _19628_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22499__B1 _21886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21514__A _21383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19559_ _23292_/Q VGND VGND VPWR VPWR _19559_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19364__B1 _19227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24353__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22570_ _22539_/X _22568_/X _20777_/X _22569_/X VGND VGND VPWR VPWR _22571_/A sky130_fd_sc_hd__o22a_4
XFILLER_55_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21521_ _21227_/A _21521_/B VGND VGND VPWR VPWR _21521_/X sky130_fd_sc_hd__or2_4
XFILLER_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18823__A _16291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24240_ _24654_/CLK _24240_/D HRESETn VGND VGND VPWR VPWR _16341_/A sky130_fd_sc_hd__dfrtp_4
X_21452_ _21452_/A VGND VGND VPWR VPWR _21452_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20403_ _20405_/A _20205_/Y VGND VGND VPWR VPWR _20403_/X sky130_fd_sc_hd__or2_4
XFILLER_135_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21383_ _21383_/A _21383_/B VGND VGND VPWR VPWR _21384_/C sky130_fd_sc_hd__or2_4
XANTENNA__22671__B1 _16073_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24171_ _24171_/CLK _24171_/D HRESETn VGND VGND VPWR VPWR _16522_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_119_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23122_ _23939_/CLK _20023_/X VGND VGND VPWR VPWR _23122_/Q sky130_fd_sc_hd__dfxtp_4
X_20334_ _20249_/A VGND VGND VPWR VPWR _20334_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16350__B1 _16087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22999__B _22999_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20265_ _23765_/Q _20265_/B VGND VGND VPWR VPWR _20266_/D sky130_fd_sc_hd__and2_4
X_23053_ _23040_/X VGND VGND VPWR VPWR IRQ[1] sky130_fd_sc_hd__buf_2
XFILLER_89_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25141__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22004_ _22004_/A _21907_/X _22004_/C _22004_/D VGND VGND VPWR VPWR HRDATA[6] sky130_fd_sc_hd__or4_4
XFILLER_62_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20196_ _20196_/A _20195_/X VGND VGND VPWR VPWR _23779_/D sky130_fd_sc_hd__or2_4
XFILLER_66_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22080__A _21519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21408__B _21408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13467__B2 _13463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23955_ _23969_/CLK _23955_/D HRESETn VGND VGND VPWR VPWR _22395_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21127__C _21123_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_9_0_HCLK clkbuf_4_4_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22906_ _22906_/A _22887_/X _22832_/C _22905_/X VGND VGND VPWR VPWR HRDATA[27] sky130_fd_sc_hd__or4_4
XFILLER_44_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12111__A _24554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23886_ _25186_/CLK _23886_/D HRESETn VGND VGND VPWR VPWR _18093_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15759__A3 _15477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22837_ _22968_/A _22837_/B VGND VGND VPWR VPWR _22851_/B sky130_fd_sc_hd__and2_4
XANTENNA__14967__B2 _24285_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16518__A _16499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22239__B _22238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15422__A _15422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24094__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13570_ _13549_/Y _13553_/X _13567_/A _13549_/A _13569_/Y VGND VGND VPWR VPWR _13570_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21162__B1 _21930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22768_ _22637_/X _22765_/Y _22601_/X _22767_/X VGND VGND VPWR VPWR _22768_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ _12509_/A _12515_/B _12520_/Y VGND VGND VPWR VPWR _12521_/X sky130_fd_sc_hd__and3_4
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24507_ _25044_/CLK _24507_/D HRESETn VGND VGND VPWR VPWR _12596_/A sky130_fd_sc_hd__dfrtp_4
X_21719_ _21719_/A VGND VGND VPWR VPWR _22226_/A sky130_fd_sc_hd__buf_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19107__B1 _19041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22699_ _22348_/X _22692_/X _22694_/X _22585_/X _22698_/Y VGND VGND VPWR VPWR _22699_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_40_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15240_ _15240_/A VGND VGND VPWR VPWR _15240_/X sky130_fd_sc_hd__buf_2
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12452_ _12434_/A _12450_/X _12451_/X VGND VGND VPWR VPWR _25095_/D sky130_fd_sc_hd__and3_4
X_24438_ _24502_/CLK _15790_/X HRESETn VGND VGND VPWR VPWR _22187_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_123_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15171_ _15105_/A _15170_/X _15147_/X VGND VGND VPWR VPWR _15171_/Y sky130_fd_sc_hd__a21oi_4
X_12383_ _12416_/A _24493_/Q _22678_/A _12382_/Y VGND VGND VPWR VPWR _12383_/X sky130_fd_sc_hd__a2bb2o_4
X_24369_ _24425_/CLK _15980_/X HRESETn VGND VGND VPWR VPWR _22192_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_125_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14122_ _14120_/B VGND VGND VPWR VPWR _14122_/X sky130_fd_sc_hd__buf_2
XFILLER_67_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14053_ _14048_/A VGND VGND VPWR VPWR _14053_/X sky130_fd_sc_hd__buf_2
X_18930_ _18929_/Y _18927_/X _18817_/X _18927_/X VGND VGND VPWR VPWR _23515_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11828__C _11694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13004_ _12925_/X _13004_/B _13003_/Y VGND VGND VPWR VPWR _13004_/X sky130_fd_sc_hd__and3_4
X_18861_ _13157_/B VGND VGND VPWR VPWR _18861_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_254_0_HCLK clkbuf_8_255_0_HCLK/A VGND VGND VPWR VPWR _24706_/CLK sky130_fd_sc_hd__clkbuf_1
X_17812_ _17944_/A _17812_/B VGND VGND VPWR VPWR _17812_/X sky130_fd_sc_hd__or2_4
X_18792_ _18792_/A VGND VGND VPWR VPWR _18792_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14955_ _14955_/A VGND VGND VPWR VPWR _15197_/A sky130_fd_sc_hd__inv_2
X_17743_ _17899_/A _17743_/B VGND VGND VPWR VPWR _17746_/B sky130_fd_sc_hd__or2_4
XFILLER_63_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12130__B2 _24559_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13906_ _24905_/Q _13892_/X _13905_/X _13825_/X _13903_/X VGND VGND VPWR VPWR _24906_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_1_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23762__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14886_ _14885_/Y _24286_/Q _14885_/Y _24286_/Q VGND VGND VPWR VPWR _14886_/X sky130_fd_sc_hd__a2bb2o_4
X_17674_ _17674_/A VGND VGND VPWR VPWR _17726_/A sky130_fd_sc_hd__inv_2
XFILLER_36_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19413_ _13313_/B VGND VGND VPWR VPWR _19413_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21334__A _21144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13837_ _13833_/A _13828_/C _13880_/C VGND VGND VPWR VPWR _13837_/X sky130_fd_sc_hd__or3_4
X_16625_ _16625_/A VGND VGND VPWR VPWR _16625_/X sky130_fd_sc_hd__buf_2
XFILLER_62_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19346__B1 _19232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22149__B _22227_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15332__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16556_ _14218_/A VGND VGND VPWR VPWR _16556_/X sky130_fd_sc_hd__buf_2
X_19344_ _19343_/Y _19341_/X _19207_/X _19341_/X VGND VGND VPWR VPWR _19344_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13768_ _13716_/C VGND VGND VPWR VPWR _13770_/B sky130_fd_sc_hd__inv_2
XFILLER_43_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19254__A2_N _19251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12719_ _12554_/X _12710_/D VGND VGND VPWR VPWR _12720_/C sky130_fd_sc_hd__nand2_4
X_15507_ HWDATA[11] VGND VGND VPWR VPWR _15507_/X sky130_fd_sc_hd__buf_2
X_16487_ _16485_/Y _16481_/X _11536_/X _16486_/X VGND VGND VPWR VPWR _16487_/X sky130_fd_sc_hd__a2bb2o_4
X_19275_ _19273_/Y _19274_/X _19227_/X _19274_/X VGND VGND VPWR VPWR _23393_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15907__B1 _15709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13699_ _13697_/X _13698_/X _14083_/A _13693_/X VGND VGND VPWR VPWR _13699_/X sky130_fd_sc_hd__o22a_4
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15438_ _15438_/A _14431_/A VGND VGND VPWR VPWR _15440_/A sky130_fd_sc_hd__or2_4
X_18226_ _18226_/A _18224_/X _18225_/Y VGND VGND VPWR VPWR _23876_/D sky130_fd_sc_hd__and3_4
XANTENNA__16580__B1 _16251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13394__B1 SCLK_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15369_ HWDATA[14] VGND VGND VPWR VPWR _15369_/X sky130_fd_sc_hd__buf_2
X_18157_ _23854_/Q VGND VGND VPWR VPWR _18312_/A sky130_fd_sc_hd__inv_2
XFILLER_8_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17259__A _17252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22653__B1 _24046_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23746__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17108_ _16992_/Y _17108_/B VGND VGND VPWR VPWR _17108_/X sky130_fd_sc_hd__or2_4
XFILLER_117_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18088_ _13049_/A _18080_/Y _18085_/X VGND VGND VPWR VPWR _23890_/D sky130_fd_sc_hd__a21oi_4
XFILLER_137_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17039_ _24041_/Q VGND VGND VPWR VPWR _17116_/A sky130_fd_sc_hd__inv_2
XFILLER_125_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20050_ _23111_/Q VGND VGND VPWR VPWR _21154_/B sky130_fd_sc_hd__inv_2
XFILLER_98_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20413__A _20413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16635__B2 _16622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15507__A HWDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24534__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23740_ _24259_/CLK _20616_/X HRESETn VGND VGND VPWR VPWR _13535_/C sky130_fd_sc_hd__dfrtp_4
X_20952_ _20946_/X _19776_/Y VGND VGND VPWR VPWR _20952_/X sky130_fd_sc_hd__or2_4
XANTENNA__16399__B1 _16141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21244__A _21396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23671_ _23680_/CLK _23671_/D HRESETn VGND VGND VPWR VPWR _23671_/Q sky130_fd_sc_hd__dfrtp_4
X_20883_ _20883_/A _15426_/X VGND VGND VPWR VPWR _20883_/X sky130_fd_sc_hd__and2_4
XPHY_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19337__B1 _19221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14792__A2_N _24099_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22622_ _24241_/Q _22147_/X _22148_/X _22621_/X VGND VGND VPWR VPWR _22622_/X sky130_fd_sc_hd__a211o_4
XPHY_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13621__B2 _13620_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11632__B1 _11631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21695__B2 _21251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22553_ _22547_/X _22550_/X _22551_/X _22552_/X VGND VGND VPWR VPWR _22554_/B sky130_fd_sc_hd__o22a_4
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21504_ _21500_/X _21503_/X _21231_/X VGND VGND VPWR VPWR _21512_/B sky130_fd_sc_hd__o21a_4
XFILLER_107_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22484_ _22484_/A _21180_/X VGND VGND VPWR VPWR _22484_/X sky130_fd_sc_hd__and2_4
XANTENNA__16571__B1 _16141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24223_ _24225_/CLK _16386_/X HRESETn VGND VGND VPWR VPWR _24223_/Q sky130_fd_sc_hd__dfrtp_4
X_21435_ _24096_/Q _21298_/B VGND VGND VPWR VPWR _21438_/B sky130_fd_sc_hd__or2_4
XANTENNA__17169__A _17086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11935__A1 _23791_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24154_ _24098_/CLK _24154_/D HRESETn VGND VGND VPWR VPWR _14814_/A sky130_fd_sc_hd__dfrtp_4
X_21366_ _21356_/Y _21365_/Y _21192_/X VGND VGND VPWR VPWR _21366_/X sky130_fd_sc_hd__o21a_4
X_23105_ _23925_/CLK _23105_/D VGND VGND VPWR VPWR _23105_/Q sky130_fd_sc_hd__dfxtp_4
X_20317_ _20317_/A VGND VGND VPWR VPWR _20317_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20670__A2 _20552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24085_ _24064_/CLK _24085_/D HRESETn VGND VGND VPWR VPWR _24085_/Q sky130_fd_sc_hd__dfrtp_4
X_21297_ _21297_/A VGND VGND VPWR VPWR _21570_/A sky130_fd_sc_hd__buf_2
X_23036_ _23036_/A _23035_/X VGND VGND VPWR VPWR _23036_/X sky130_fd_sc_hd__and2_4
X_20248_ _20244_/X _20247_/X VGND VGND VPWR VPWR _23769_/D sky130_fd_sc_hd__or2_4
XFILLER_77_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16626__B2 _16622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15417__A _14197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11945__A _11944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20179_ _23777_/Q _20179_/B _20179_/C _20249_/B VGND VGND VPWR VPWR _20179_/X sky130_fd_sc_hd__and4_4
XFILLER_114_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_8_0_HCLK_A clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_21_0_HCLK clkbuf_8_21_0_HCLK/A VGND VGND VPWR VPWR _24824_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22850__A1_N _21546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24987_ _24953_/CLK _24987_/D HRESETn VGND VGND VPWR VPWR _24987_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21907__C1 _21895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_84_0_HCLK clkbuf_8_85_0_HCLK/A VGND VGND VPWR VPWR _24769_/CLK sky130_fd_sc_hd__clkbuf_1
X_14740_ _14740_/A VGND VGND VPWR VPWR _14740_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24275__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11952_ _11950_/X _16038_/B _22510_/B VGND VGND VPWR VPWR _11952_/X sky130_fd_sc_hd__or3_4
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23938_ _23343_/CLK _17652_/X HRESETn VGND VGND VPWR VPWR _23938_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24204__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14671_ _14671_/A VGND VGND VPWR VPWR _14671_/Y sky130_fd_sc_hd__inv_2
X_11883_ _11883_/A _11894_/A VGND VGND VPWR VPWR _11884_/B sky130_fd_sc_hd__and2_4
XANTENNA__23898__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23869_ _23872_/CLK _23869_/D HRESETn VGND VGND VPWR VPWR _23869_/Q sky130_fd_sc_hd__dfrtp_4
X_16410_ _16408_/Y _16409_/X _16153_/X _16409_/X VGND VGND VPWR VPWR _16410_/X sky130_fd_sc_hd__a2bb2o_4
X_13622_ _13622_/A VGND VGND VPWR VPWR _13622_/Y sky130_fd_sc_hd__inv_2
X_17390_ _17390_/A _17386_/X _17389_/Y VGND VGND VPWR VPWR _17390_/X sky130_fd_sc_hd__and3_4
XFILLER_38_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16341_ _16341_/A VGND VGND VPWR VPWR _16341_/Y sky130_fd_sc_hd__inv_2
X_13553_ _13580_/A VGND VGND VPWR VPWR _13553_/X sky130_fd_sc_hd__buf_2
X_12504_ _12403_/B _12503_/X VGND VGND VPWR VPWR _12505_/B sky130_fd_sc_hd__or2_4
X_19060_ _19055_/Y _19058_/X _19059_/X _19058_/X VGND VGND VPWR VPWR _23470_/D sky130_fd_sc_hd__a2bb2o_4
X_16272_ _16268_/X _16269_/X _16087_/A _22477_/A _16270_/X VGND VGND VPWR VPWR _16272_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_16_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13484_ _13468_/A _13468_/B VGND VGND VPWR VPWR _13484_/X sky130_fd_sc_hd__or2_4
XFILLER_125_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15223_ _15110_/B _15222_/X VGND VGND VPWR VPWR _15224_/B sky130_fd_sc_hd__or2_4
X_18011_ _18011_/A VGND VGND VPWR VPWR _18011_/Y sky130_fd_sc_hd__inv_2
X_12435_ _12401_/B _12424_/X _12427_/X _12432_/B VGND VGND VPWR VPWR _12435_/X sky130_fd_sc_hd__a211o_4
XFILLER_16_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25063__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15154_ _15154_/A _15154_/B _15153_/X VGND VGND VPWR VPWR _24673_/D sky130_fd_sc_hd__and3_4
X_12366_ _12497_/A VGND VGND VPWR VPWR _12413_/A sky130_fd_sc_hd__inv_2
XFILLER_114_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14105_ _23126_/Q _14100_/X _14104_/A _23655_/D _14104_/Y VGND VGND VPWR VPWR _24854_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_113_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15085_ _15085_/A _15123_/B VGND VGND VPWR VPWR _15085_/X sky130_fd_sc_hd__or2_4
X_19962_ _23144_/Q VGND VGND VPWR VPWR _19962_/Y sky130_fd_sc_hd__inv_2
X_12297_ _12293_/B _12297_/B _12300_/C VGND VGND VPWR VPWR _12297_/X sky130_fd_sc_hd__and3_4
X_14036_ _24875_/Q VGND VGND VPWR VPWR _14036_/Y sky130_fd_sc_hd__inv_2
X_18913_ _18899_/Y VGND VGND VPWR VPWR _18913_/X sky130_fd_sc_hd__buf_2
XANTENNA__21329__A _21333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19893_ _21673_/B _19890_/X _19825_/X _19890_/X VGND VGND VPWR VPWR _23171_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18844_ _23545_/Q VGND VGND VPWR VPWR _21375_/B sky130_fd_sc_hd__inv_2
XFILLER_121_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14231__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18775_ _23569_/Q VGND VGND VPWR VPWR _18775_/Y sky130_fd_sc_hd__inv_2
X_15987_ _15987_/A VGND VGND VPWR VPWR _15987_/X sky130_fd_sc_hd__buf_2
XANTENNA__22166__A2 _22488_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20887__B _20931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17726_ _17726_/A VGND VGND VPWR VPWR _17780_/A sky130_fd_sc_hd__buf_2
XANTENNA__17542__A _17481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14938_ _24651_/Q _14936_/Y _15218_/A _14937_/Y VGND VGND VPWR VPWR _14943_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21064__A _15821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17657_ _13407_/B VGND VGND VPWR VPWR _17657_/Y sky130_fd_sc_hd__inv_2
X_14869_ _14869_/A _14869_/B VGND VGND VPWR VPWR _14873_/B sky130_fd_sc_hd__or2_4
XANTENNA__16158__A _16165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11590__A _16093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16608_ _16608_/A VGND VGND VPWR VPWR _16608_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21999__A _16685_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17588_ _21839_/A _17587_/X VGND VGND VPWR VPWR _17594_/B sky130_fd_sc_hd__or2_4
XFILLER_95_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23998__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19327_ _19327_/A VGND VGND VPWR VPWR _19327_/Y sky130_fd_sc_hd__inv_2
X_16539_ _16539_/A VGND VGND VPWR VPWR _16539_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23927__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19258_ _22047_/A VGND VGND VPWR VPWR _19258_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13367__B1 _11612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18209_ _18209_/A VGND VGND VPWR VPWR _18218_/B sky130_fd_sc_hd__inv_2
X_19189_ _19144_/A _19189_/B _19100_/A VGND VGND VPWR VPWR _19189_/X sky130_fd_sc_hd__or3_4
XANTENNA__13310__A _13102_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21220_ _14443_/B VGND VGND VPWR VPWR _21385_/A sky130_fd_sc_hd__buf_2
XANTENNA__20101__B2 _20098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21151_ _17629_/B VGND VGND VPWR VPWR _21340_/A sky130_fd_sc_hd__buf_2
XANTENNA__16043__D _22265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16621__A _16621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22929__A1 _16054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20102_ _23091_/Q VGND VGND VPWR VPWR _20102_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21082_ _24874_/Q _21082_/B VGND VGND VPWR VPWR _21082_/X sky130_fd_sc_hd__and2_4
XANTENNA__24786__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20033_ _20033_/A VGND VGND VPWR VPWR _22107_/B sky130_fd_sc_hd__inv_2
X_24910_ _24904_/CLK _24910_/D HRESETn VGND VGND VPWR VPWR _13827_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24715__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_1_0_HCLK_A clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24841_ _24841_/CLK _24841_/D HRESETn VGND VGND VPWR VPWR _24841_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15292__B1 _15291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19558__B1 _11839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24772_ _24776_/CLK _24772_/D HRESETn VGND VGND VPWR VPWR _24772_/Q sky130_fd_sc_hd__dfrtp_4
X_21984_ _22036_/A VGND VGND VPWR VPWR _21984_/X sky130_fd_sc_hd__buf_2
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23723_ _24606_/CLK _23723_/D HRESETn VGND VGND VPWR VPWR _20542_/B sky130_fd_sc_hd__dfrtp_4
X_20935_ _20935_/A VGND VGND VPWR VPWR _20935_/Y sky130_fd_sc_hd__inv_2
XPHY_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12596__A _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23654_ _24879_/CLK _23654_/D HRESETn VGND VGND VPWR VPWR _23654_/Q sky130_fd_sc_hd__dfrtp_4
X_20866_ _20866_/A VGND VGND VPWR VPWR _20866_/X sky130_fd_sc_hd__buf_2
XPHY_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22605_ _22605_/A _22527_/B VGND VGND VPWR VPWR _22605_/X sky130_fd_sc_hd__and2_4
XANTENNA__11605__B1 _11604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23668__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23585_ _23586_/CLK _23585_/D VGND VGND VPWR VPWR _17888_/B sky130_fd_sc_hd__dfxtp_4
X_20797_ _21285_/B VGND VGND VPWR VPWR _22870_/B sky130_fd_sc_hd__buf_2
XPHY_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22536_ _21972_/X VGND VGND VPWR VPWR _22536_/X sky130_fd_sc_hd__buf_2
XFILLER_126_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22467_ _21042_/X _22466_/X _22197_/X _24410_/Q _21047_/X VGND VGND VPWR VPWR _22468_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_10_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12220_ _12190_/A _12216_/X _12219_/Y VGND VGND VPWR VPWR _25126_/D sky130_fd_sc_hd__and3_4
X_24206_ _24244_/CLK _24206_/D HRESETn VGND VGND VPWR VPWR _24206_/Q sky130_fd_sc_hd__dfrtp_4
X_21418_ _21432_/A VGND VGND VPWR VPWR _22155_/A sky130_fd_sc_hd__buf_2
X_25186_ _25186_/CLK _11768_/Y HRESETn VGND VGND VPWR VPWR _11716_/A sky130_fd_sc_hd__dfstp_4
X_22398_ _21246_/X _22395_/X _22398_/C _22398_/D VGND VGND VPWR VPWR _22398_/X sky130_fd_sc_hd__or4_4
XFILLER_135_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12151_ _12142_/X _12151_/B _12147_/X _12150_/X VGND VGND VPWR VPWR _12161_/C sky130_fd_sc_hd__or4_4
X_24137_ _24094_/CLK _16600_/X HRESETn VGND VGND VPWR VPWR _24137_/Q sky130_fd_sc_hd__dfrtp_4
X_21349_ _21935_/A _21349_/B VGND VGND VPWR VPWR _21349_/X sky130_fd_sc_hd__or2_4
XANTENNA__19729__A2_N _19727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21149__A _21339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12082_ _12082_/A VGND VGND VPWR VPWR _12083_/A sky130_fd_sc_hd__inv_2
XFILLER_78_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24068_ _24620_/CLK _16934_/X HRESETn VGND VGND VPWR VPWR _16776_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_49_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12333__B2 _12332_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15910_ _15916_/A _16127_/A VGND VGND VPWR VPWR _15910_/X sky130_fd_sc_hd__or2_4
XANTENNA__24456__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23019_ _22334_/A _23019_/B _23019_/C VGND VGND VPWR VPWR _23030_/B sky130_fd_sc_hd__and3_4
X_16890_ _16890_/A _16888_/X _16889_/X VGND VGND VPWR VPWR _24080_/D sky130_fd_sc_hd__and3_4
X_15841_ _24421_/Q VGND VGND VPWR VPWR _15841_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15283__B1 _15282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18560_ _18484_/A _18551_/B _18559_/X VGND VGND VPWR VPWR _18560_/X sky130_fd_sc_hd__and3_4
XANTENNA__20159__A1 _24822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12984_ _12984_/A _12984_/B VGND VGND VPWR VPWR _12984_/X sky130_fd_sc_hd__or2_4
X_15772_ HWDATA[19] VGND VGND VPWR VPWR _15772_/X sky130_fd_sc_hd__buf_2
XANTENNA__21356__B1 _21175_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22174__A1_N _16700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17511_ _17505_/D _17511_/B VGND VGND VPWR VPWR _17511_/X sky130_fd_sc_hd__or2_4
X_11935_ _23791_/Q _11918_/A _20880_/A _11931_/X VGND VGND VPWR VPWR _11935_/X sky130_fd_sc_hd__o22a_4
X_14723_ _24700_/Q _14722_/A _15035_/A _14722_/Y VGND VGND VPWR VPWR _14734_/A sky130_fd_sc_hd__o22a_4
XFILLER_73_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18491_ _18491_/A _18491_/B VGND VGND VPWR VPWR _18492_/C sky130_fd_sc_hd__or2_4
XFILLER_17_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14654_ _14621_/X _14653_/X _15284_/A _14647_/X VGND VGND VPWR VPWR _14654_/Y sky130_fd_sc_hd__a22oi_4
X_17442_ _23979_/Q _17441_/Y VGND VGND VPWR VPWR _17443_/B sky130_fd_sc_hd__or2_4
X_11866_ _11871_/C _11871_/D VGND VGND VPWR VPWR _11866_/X sky130_fd_sc_hd__and2_4
XANTENNA__21108__B1 _21107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13605_ _13555_/B _13604_/X _13553_/X _13586_/X _11676_/A VGND VGND VPWR VPWR _24948_/D
+ sky130_fd_sc_hd__a32o_4
X_14585_ _24732_/Q VGND VGND VPWR VPWR _14587_/A sky130_fd_sc_hd__inv_2
X_17373_ _17286_/Y _17373_/B VGND VGND VPWR VPWR _17373_/X sky130_fd_sc_hd__or2_4
X_11797_ _11797_/A VGND VGND VPWR VPWR _11797_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18193__A _18485_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19112_ _19111_/Y _19106_/X _19089_/X _19106_/X VGND VGND VPWR VPWR _19112_/X sky130_fd_sc_hd__a2bb2o_4
X_13536_ _23742_/Q _20617_/A _13535_/X VGND VGND VPWR VPWR _13537_/C sky130_fd_sc_hd__or3_4
X_16324_ _16323_/Y _16321_/X _15479_/X _16321_/X VGND VGND VPWR VPWR _16324_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13349__B1 _11631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16255_ _14960_/Y _16247_/X _16254_/X _16247_/X VGND VGND VPWR VPWR _16255_/X sky130_fd_sc_hd__a2bb2o_4
X_19043_ _19040_/Y _19035_/X _19041_/X _19042_/X VGND VGND VPWR VPWR _19043_/X sky130_fd_sc_hd__a2bb2o_4
X_13467_ _13465_/Y _13463_/Y _21696_/A _13463_/A VGND VGND VPWR VPWR _13468_/B sky130_fd_sc_hd__o22a_4
X_15206_ _15109_/Y _15203_/B VGND VGND VPWR VPWR _15207_/C sky130_fd_sc_hd__nand2_4
X_12418_ _12391_/Y _12401_/X _12418_/C _12424_/A VGND VGND VPWR VPWR _12419_/A sky130_fd_sc_hd__or4_4
X_16186_ _16186_/A VGND VGND VPWR VPWR _16186_/Y sky130_fd_sc_hd__inv_2
X_13398_ _13398_/A VGND VGND VPWR VPWR _13398_/X sky130_fd_sc_hd__buf_2
XFILLER_86_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15137_ _14946_/Y _15152_/A VGND VGND VPWR VPWR _15154_/B sky130_fd_sc_hd__or2_4
X_12349_ _12349_/A VGND VGND VPWR VPWR _12349_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15068_ _14839_/Y _15067_/X _15027_/X _15063_/B VGND VGND VPWR VPWR _15068_/X sky130_fd_sc_hd__a211o_4
X_19945_ _23150_/Q VGND VGND VPWR VPWR _19945_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21059__A _22933_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14019_ _24622_/Q _15314_/B VGND VGND VPWR VPWR _16038_/D sky130_fd_sc_hd__or2_4
XANTENNA__11585__A _11585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24197__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19876_ _19876_/A VGND VGND VPWR VPWR _19876_/X sky130_fd_sc_hd__buf_2
XFILLER_95_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17263__A1 _25199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24126__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18827_ _18827_/A VGND VGND VPWR VPWR _18827_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15274__B1 _14232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22139__A2 _22011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18758_ _17671_/B VGND VGND VPWR VPWR _18758_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21347__B1 _21930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17709_ _14563_/A VGND VGND VPWR VPWR _17815_/A sky130_fd_sc_hd__buf_2
XANTENNA__17015__B2 _17027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18689_ _23598_/Q VGND VGND VPWR VPWR _18689_/Y sky130_fd_sc_hd__inv_2
X_20720_ _20720_/A VGND VGND VPWR VPWR _20720_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21522__A _21235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20651_ _20651_/A VGND VGND VPWR VPWR _20651_/X sky130_fd_sc_hd__buf_2
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23761__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16616__A _24126_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15520__A _11625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23370_ _23374_/CLK _19339_/X VGND VGND VPWR VPWR _23370_/Q sky130_fd_sc_hd__dfxtp_4
X_20582_ _20582_/A VGND VGND VPWR VPWR _20582_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16526__B1 _16096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11602__A3 _15788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22321_ _22354_/A _22320_/X VGND VGND VPWR VPWR _22321_/Y sky130_fd_sc_hd__nor2_4
XFILLER_104_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25040_ _25044_/CLK _12766_/X HRESETn VGND VGND VPWR VPWR _25040_/Q sky130_fd_sc_hd__dfrtp_4
X_22252_ _15463_/X _22250_/X _22251_/X _24555_/Q _15824_/A VGND VGND VPWR VPWR _22252_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12012__B1 _11643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24967__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18550__B _18468_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21203_ _21238_/A VGND VGND VPWR VPWR _21374_/A sky130_fd_sc_hd__buf_2
XFILLER_69_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17447__A _17446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22183_ _22183_/A _22183_/B _22168_/X _22182_/X VGND VGND VPWR VPWR HRDATA[8] sky130_fd_sc_hd__or4_4
X_21134_ _21352_/A _21134_/B VGND VGND VPWR VPWR _21134_/X sky130_fd_sc_hd__or2_4
XFILLER_59_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21065_ _21064_/Y VGND VGND VPWR VPWR _21066_/B sky130_fd_sc_hd__buf_2
XFILLER_8_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20016_ _22092_/B _20015_/X _19711_/X _20015_/X VGND VGND VPWR VPWR _20016_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24824_ _24824_/CLK _14192_/X HRESETn VGND VGND VPWR VPWR _24824_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21338__B1 _17639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14715__A1_N _14712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24755_ _24757_/CLK _24755_/D HRESETn VGND VGND VPWR VPWR _13447_/A sky130_fd_sc_hd__dfrtp_4
X_21967_ _21967_/A VGND VGND VPWR VPWR _21967_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23849__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _24622_/Q _11951_/B _14020_/A VGND VGND VPWR VPWR _11720_/X sky130_fd_sc_hd__or3_4
XANTENNA__22550__A2 _22537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19951__B1 _19421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23706_ _23706_/CLK _20471_/X HRESETn VGND VGND VPWR VPWR _20468_/A sky130_fd_sc_hd__dfrtp_4
X_20918_ _20917_/X VGND VGND VPWR VPWR _20918_/X sky130_fd_sc_hd__buf_2
XFILLER_42_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24686_ _24674_/CLK _24686_/D HRESETn VGND VGND VPWR VPWR _24686_/Q sky130_fd_sc_hd__dfrtp_4
X_21898_ _21898_/A _21106_/X VGND VGND VPWR VPWR _21898_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_158_0_HCLK clkbuf_7_79_0_HCLK/X VGND VGND VPWR VPWR _24451_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _24958_/Q VGND VGND VPWR VPWR _13564_/A sky130_fd_sc_hd__inv_2
XFILLER_70_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23637_ _24811_/CLK _20313_/Y HRESETn VGND VGND VPWR VPWR _18615_/A sky130_fd_sc_hd__dfrtp_4
X_20849_ _20849_/A _20849_/B _20846_/X _20849_/D VGND VGND VPWR VPWR _20850_/A sky130_fd_sc_hd__or4_4
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15430__A _15430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14370_ _14369_/X VGND VGND VPWR VPWR _14390_/D sky130_fd_sc_hd__inv_2
XFILLER_11_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11582_ _11579_/Y _11577_/X _11581_/X _11577_/X VGND VGND VPWR VPWR _11582_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23568_ _23568_/CLK _18779_/X VGND VGND VPWR VPWR _17924_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13321_ _13057_/A _13320_/X _24996_/Q _13054_/X VGND VGND VPWR VPWR _24996_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19259__D _22024_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23666__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22519_ _22364_/X _22518_/X _21981_/X _24518_/Q _22366_/X VGND VGND VPWR VPWR _22519_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24752__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23499_ _23586_/CLK _18978_/X VGND VGND VPWR VPWR _13161_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_7_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16040_ _21882_/A VGND VGND VPWR VPWR _21273_/A sky130_fd_sc_hd__inv_2
XFILLER_100_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13252_ _13110_/A _23321_/Q VGND VGND VPWR VPWR _13253_/C sky130_fd_sc_hd__or2_4
XFILLER_129_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12003__B1 _11626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22263__A _22223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12203_ _12538_/B VGND VGND VPWR VPWR _12203_/X sky130_fd_sc_hd__buf_2
X_13183_ _13146_/A _19404_/A VGND VGND VPWR VPWR _13183_/X sky130_fd_sc_hd__or2_4
XANTENNA__24637__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25169_ _23288_/CLK _25169_/D HRESETn VGND VGND VPWR VPWR _25169_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16261__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12134_ _25125_/Q VGND VGND VPWR VPWR _12207_/A sky130_fd_sc_hd__inv_2
X_17991_ _17982_/X _17990_/X _16451_/X _22215_/A _17983_/X VGND VGND VPWR VPWR _17991_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_78_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19730_ _19730_/A VGND VGND VPWR VPWR _21132_/B sky130_fd_sc_hd__inv_2
XANTENNA__24290__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12065_ _12065_/A VGND VGND VPWR VPWR _16559_/A sky130_fd_sc_hd__buf_2
X_16942_ _16942_/A VGND VGND VPWR VPWR _16942_/Y sky130_fd_sc_hd__inv_2
X_19661_ _19661_/A VGND VGND VPWR VPWR _19661_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16873_ _16863_/A _16875_/B _16872_/Y VGND VGND VPWR VPWR _16873_/X sky130_fd_sc_hd__o21a_4
XFILLER_133_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20511__A _20511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18612_ _20297_/A _20293_/A VGND VGND VPWR VPWR _20298_/A sky130_fd_sc_hd__or2_4
X_15824_ _15824_/A _16135_/B VGND VGND VPWR VPWR _15824_/X sky130_fd_sc_hd__and2_4
X_19592_ _19592_/A VGND VGND VPWR VPWR _21013_/B sky130_fd_sc_hd__inv_2
XFILLER_37_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18543_ _18543_/A _18543_/B VGND VGND VPWR VPWR _18544_/C sky130_fd_sc_hd__nand2_4
Xclkbuf_7_54_0_HCLK clkbuf_7_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_54_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12967_ _12836_/Y _12964_/X VGND VGND VPWR VPWR _12967_/X sky130_fd_sc_hd__or2_4
X_15755_ _12849_/Y _15752_/X _15332_/X _15752_/X VGND VGND VPWR VPWR _15755_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20001__B1 _15522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19942__B1 _15561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13125__A _13065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11918_ _11918_/A VGND VGND VPWR VPWR _11919_/A sky130_fd_sc_hd__inv_2
X_14706_ _24698_/Q VGND VGND VPWR VPWR _14876_/D sky130_fd_sc_hd__inv_2
XANTENNA__17820__A _17721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18474_ _18463_/A _18474_/B _18473_/X VGND VGND VPWR VPWR _23838_/D sky130_fd_sc_hd__and3_4
X_12898_ _12898_/A VGND VGND VPWR VPWR _12898_/Y sky130_fd_sc_hd__inv_2
X_15686_ _15684_/X _15672_/X _15494_/X _24483_/Q _15685_/X VGND VGND VPWR VPWR _24483_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_61_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22438__A _22438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17425_ _17423_/A _17413_/B _17425_/C VGND VGND VPWR VPWR _17425_/X sky130_fd_sc_hd__and3_4
XANTENNA__21342__A _21342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11849_ _11847_/Y _11840_/X _11848_/X _11840_/X VGND VGND VPWR VPWR _11849_/X sky130_fd_sc_hd__a2bb2o_4
X_14637_ _14620_/A VGND VGND VPWR VPWR _14643_/A sky130_fd_sc_hd__buf_2
XFILLER_57_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14568_ _17732_/A VGND VGND VPWR VPWR _14569_/A sky130_fd_sc_hd__buf_2
X_17356_ _17622_/B _17352_/B _17355_/X VGND VGND VPWR VPWR _17356_/X sky130_fd_sc_hd__or3_4
XFILLER_105_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20304__A1 _14264_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16307_ _16313_/A VGND VGND VPWR VPWR _16308_/A sky130_fd_sc_hd__buf_2
X_13519_ _13519_/A VGND VGND VPWR VPWR _13519_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13990__B1 _24812_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14499_ _14498_/X VGND VGND VPWR VPWR _24751_/D sky130_fd_sc_hd__inv_2
X_17287_ _11544_/Y _24004_/Q _11562_/A _17286_/Y VGND VGND VPWR VPWR _17290_/C sky130_fd_sc_hd__a2bb2o_4
X_19026_ _21374_/B _19025_/X _15563_/X _19025_/X VGND VGND VPWR VPWR _23481_/D sky130_fd_sc_hd__a2bb2o_4
X_16238_ _16228_/X _16234_/X _15743_/X _24286_/Q _16237_/X VGND VGND VPWR VPWR _24286_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_127_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22173__A _21069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20068__B1 _19808_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12545__B2 _24533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24378__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16169_ _24308_/Q VGND VGND VPWR VPWR _16169_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23006__B1 _24533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24307__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19928_ _22064_/B _19927_/X _19442_/A _19927_/X VGND VGND VPWR VPWR _23158_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21568__B1 _21107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19859_ _19859_/A VGND VGND VPWR VPWR _19859_/X sky130_fd_sc_hd__buf_2
XFILLER_110_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22780__A2 _20799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22870_ _15337_/Y _22870_/B VGND VGND VPWR VPWR _22870_/X sky130_fd_sc_hd__and2_4
XANTENNA__20791__A1 _21448_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20791__B2 _11940_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21821_ _21817_/X _21820_/X _20968_/X VGND VGND VPWR VPWR _21821_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_83_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23942__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19933__B1 _19448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25166__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24540_ _23179_/CLK _24540_/D HRESETn VGND VGND VPWR VPWR _19818_/A sky130_fd_sc_hd__dfrtp_4
X_21752_ _21752_/A _19279_/Y _21752_/C VGND VGND VPWR VPWR _21752_/X sky130_fd_sc_hd__and3_4
XFILLER_58_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22348__A _23023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21740__B1 _24805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20703_ scl_oen_o_S4 _20703_/B VGND VGND VPWR VPWR _20703_/X sky130_fd_sc_hd__and2_4
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24471_ _24307_/CLK _24471_/D HRESETn VGND VGND VPWR VPWR _21567_/A sky130_fd_sc_hd__dfrtp_4
X_21683_ _21667_/X _21683_/B VGND VGND VPWR VPWR _21683_/X sky130_fd_sc_hd__or2_4
XFILLER_51_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23422_ _23596_/CLK _19192_/X VGND VGND VPWR VPWR _23422_/Q sky130_fd_sc_hd__dfxtp_4
X_20634_ _20635_/B VGND VGND VPWR VPWR _20634_/Y sky130_fd_sc_hd__inv_2
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23353_ _23353_/CLK _19388_/X VGND VGND VPWR VPWR _19385_/A sky130_fd_sc_hd__dfxtp_4
X_20565_ _20564_/X VGND VGND VPWR VPWR _23729_/D sky130_fd_sc_hd__inv_2
XFILLER_137_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18561__A pwm_S7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22304_ _13360_/A _22303_/X _22251_/X _24556_/Q _15824_/A VGND VGND VPWR VPWR _22304_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22048__B2 _21400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23284_ _23308_/CLK _19582_/X VGND VGND VPWR VPWR _23284_/Q sky130_fd_sc_hd__dfxtp_4
X_20496_ _20499_/A _20491_/X _20495_/X VGND VGND VPWR VPWR _20496_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__22083__A _11532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16097__A2_N _16090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25023_ _24445_/CLK _12949_/X HRESETn VGND VGND VPWR VPWR _22605_/A sky130_fd_sc_hd__dfrtp_4
X_22235_ _22730_/A _22235_/B VGND VGND VPWR VPWR _22235_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24730__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24048__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22166_ _24403_/Q _22488_/B _20782_/A _22165_/X VGND VGND VPWR VPWR _22167_/C sky130_fd_sc_hd__a211o_4
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15486__B1 _11558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21117_ _13324_/X _21116_/X VGND VGND VPWR VPWR _21117_/X sky130_fd_sc_hd__or2_4
XFILLER_117_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19392__A _15431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22097_ _17639_/A _22093_/X _22096_/X VGND VGND VPWR VPWR _22097_/X sky130_fd_sc_hd__or3_4
XFILLER_82_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12114__A _24547_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21023__A2 _21018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21048_ _21042_/X _21044_/X _21046_/X _25191_/Q _21047_/X VGND VGND VPWR VPWR _21049_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22220__B2 _21870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20331__A _20331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11953__A _11952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13870_ _13870_/A VGND VGND VPWR VPWR _14357_/B sky130_fd_sc_hd__inv_2
XANTENNA__23064__D scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12821_ _12811_/X _12821_/B _12821_/C _12821_/D VGND VGND VPWR VPWR _12821_/X sky130_fd_sc_hd__or4_4
XFILLER_90_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24807_ _23774_/CLK _14250_/X HRESETn VGND VGND VPWR VPWR _14247_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__23683__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22999_ _22999_/A _22999_/B VGND VGND VPWR VPWR _22999_/X sky130_fd_sc_hd__or2_4
X_12752_ _12647_/C _12739_/X VGND VGND VPWR VPWR _12753_/C sky130_fd_sc_hd__nand2_4
X_15540_ _19445_/A VGND VGND VPWR VPWR _15540_/Y sky130_fd_sc_hd__inv_2
XPHY_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24738_ _23469_/CLK _14562_/X HRESETn VGND VGND VPWR VPWR _17806_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22258__A _22258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _18638_/B _11702_/X VGND VGND VPWR VPWR _11703_/X sky130_fd_sc_hd__or2_4
XFILLER_72_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _15470_/Y VGND VGND VPWR VPWR _15472_/A sky130_fd_sc_hd__buf_2
X_12683_ _12637_/X _12683_/B _12683_/C VGND VGND VPWR VPWR _25064_/D sky130_fd_sc_hd__and3_4
XPHY_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24669_ _24671_/CLK _24669_/D HRESETn VGND VGND VPWR VPWR _24669_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _14374_/A _14373_/Y VGND VGND VPWR VPWR _14422_/Y sky130_fd_sc_hd__nand2_4
X_17210_ _24015_/Q VGND VGND VPWR VPWR _17210_/Y sky130_fd_sc_hd__inv_2
XPHY_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ HWDATA[2] VGND VGND VPWR VPWR _11635_/A sky130_fd_sc_hd__buf_2
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18190_ _18190_/A _18190_/B _18190_/C _18189_/X VGND VGND VPWR VPWR _18190_/X sky130_fd_sc_hd__or4_4
XFILLER_30_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24889__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14353_ _14353_/A VGND VGND VPWR VPWR _14353_/Y sky130_fd_sc_hd__inv_2
X_17141_ _17034_/A _17145_/A _17144_/A _17153_/B VGND VGND VPWR VPWR _17141_/X sky130_fd_sc_hd__or4_4
XANTENNA__12775__B2 _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11565_ _11565_/A VGND VGND VPWR VPWR _11565_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24818__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13304_ _13155_/X _13304_/B _13304_/C VGND VGND VPWR VPWR _13304_/X sky130_fd_sc_hd__and3_4
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17072_ _17056_/Y VGND VGND VPWR VPWR _17074_/A sky130_fd_sc_hd__buf_2
X_14284_ _24792_/Q VGND VGND VPWR VPWR _14284_/Y sky130_fd_sc_hd__inv_2
X_11496_ _11496_/A VGND VGND VPWR VPWR _11496_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13235_ _13203_/A _13235_/B _13235_/C VGND VGND VPWR VPWR _13239_/B sky130_fd_sc_hd__and3_4
X_16023_ _17806_/A _14581_/A _16022_/Y _14581_/Y VGND VGND VPWR VPWR _16023_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17087__A _17086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24471__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21798__B1 _21868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24400__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13166_ _13166_/A _23595_/Q VGND VGND VPWR VPWR _13166_/X sky130_fd_sc_hd__or2_4
XANTENNA__18663__B1 _18662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20065__A3 _18000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12117_ _12117_/A VGND VGND VPWR VPWR _12117_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13097_ _13244_/A _13097_/B VGND VGND VPWR VPWR _13097_/X sky130_fd_sc_hd__or2_4
X_17974_ _17973_/X _12065_/A VGND VGND VPWR VPWR _17974_/X sky130_fd_sc_hd__or2_4
XANTENNA__22440__B _22859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19713_ _19713_/A VGND VGND VPWR VPWR _21916_/B sky130_fd_sc_hd__inv_2
X_12048_ _12048_/A _12048_/B _18111_/C _24835_/Q VGND VGND VPWR VPWR _12048_/X sky130_fd_sc_hd__and4_4
X_16925_ _16771_/Y _16937_/B VGND VGND VPWR VPWR _16938_/B sky130_fd_sc_hd__or2_4
XFILLER_133_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19644_ _18023_/X VGND VGND VPWR VPWR _19644_/X sky130_fd_sc_hd__buf_2
X_16856_ _16774_/Y _16854_/A VGND VGND VPWR VPWR _16856_/X sky130_fd_sc_hd__or2_4
XFILLER_20_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15807_ _15807_/A _15713_/A VGND VGND VPWR VPWR _15807_/X sky130_fd_sc_hd__or2_4
X_19575_ _19575_/A VGND VGND VPWR VPWR _19575_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16787_ _24064_/Q VGND VGND VPWR VPWR _16923_/A sky130_fd_sc_hd__inv_2
XFILLER_94_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13999_ _13999_/A VGND VGND VPWR VPWR _14000_/B sky130_fd_sc_hd__buf_2
XFILLER_46_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18526_ _18426_/X _18543_/B VGND VGND VPWR VPWR _18529_/B sky130_fd_sc_hd__or2_4
XFILLER_80_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15738_ _15418_/A _15741_/B VGND VGND VPWR VPWR _15738_/X sky130_fd_sc_hd__or2_4
XFILLER_61_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21072__A _21072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18457_ _18452_/C _18446_/X _18449_/X _18453_/Y VGND VGND VPWR VPWR _18458_/A sky130_fd_sc_hd__a211o_4
X_15669_ _15666_/A VGND VGND VPWR VPWR _15669_/X sky130_fd_sc_hd__buf_2
XFILLER_33_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_141_0_HCLK clkbuf_7_70_0_HCLK/X VGND VGND VPWR VPWR _25067_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_21_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17408_ _17320_/A _17264_/Y _17323_/C _17408_/D VGND VGND VPWR VPWR _17409_/B sky130_fd_sc_hd__or4_4
XANTENNA__21074__A2_N _13333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18388_ _18388_/A VGND VGND VPWR VPWR _18479_/A sky130_fd_sc_hd__buf_2
X_17339_ _17329_/A _17328_/X VGND VGND VPWR VPWR _17339_/X sky130_fd_sc_hd__or2_4
XANTENNA__20828__A2 _20826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24559__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22615__B _22574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20350_ _17173_/B _20350_/B _20349_/X VGND VGND VPWR VPWR _20350_/X sky130_fd_sc_hd__and3_4
XANTENNA__20416__A _20416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21089__A2_N _21043_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19009_ _23486_/Q VGND VGND VPWR VPWR _19009_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20281_ _20281_/A VGND VGND VPWR VPWR _23630_/D sky130_fd_sc_hd__inv_2
XFILLER_66_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11526__A2_N _11521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22020_ _21882_/X _22016_/X _22017_/X _22019_/X VGND VGND VPWR VPWR _22020_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20056__A3 _13663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24141__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17725__A _17725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23971_ _24361_/CLK _23971_/D HRESETn VGND VGND VPWR VPWR _16710_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_130_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13494__A2 _13492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22922_ _12401_/B _22259_/X _24055_/Q _22433_/A VGND VGND VPWR VPWR _22923_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20764__A1 _22014_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20764__B2 _21591_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22853_ _22853_/A _23004_/A VGND VGND VPWR VPWR _22853_/X sky130_fd_sc_hd__and2_4
XANTENNA__18556__A _18484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21804_ _17451_/Y _23104_/Q _21805_/A _20064_/X VGND VGND VPWR VPWR _21804_/X sky130_fd_sc_hd__o22a_4
X_22784_ _25214_/Q _20821_/X _20801_/X _22783_/X VGND VGND VPWR VPWR _22784_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21713__B1 _21175_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24523_ _24523_/CLK _24523_/D HRESETn VGND VGND VPWR VPWR _24523_/Q sky130_fd_sc_hd__dfrtp_4
X_21735_ _17204_/Y _22439_/B _23654_/Q _21088_/X VGND VGND VPWR VPWR _21737_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24454_ _24459_/CLK _15760_/X HRESETn VGND VGND VPWR VPWR _24454_/Q sky130_fd_sc_hd__dfrtp_4
X_21666_ _21010_/A VGND VGND VPWR VPWR _21675_/A sky130_fd_sc_hd__buf_2
XANTENNA__24982__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23405_ _23383_/CLK _19242_/X VGND VGND VPWR VPWR _19241_/A sky130_fd_sc_hd__dfxtp_4
X_20617_ _20617_/A VGND VGND VPWR VPWR _20617_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19387__A _11635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24911__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24385_ _24385_/CLK _15939_/X HRESETn VGND VGND VPWR VPWR _22820_/A sky130_fd_sc_hd__dfrtp_4
X_21597_ _12972_/A _15576_/X _23946_/Q _21990_/A VGND VGND VPWR VPWR _21597_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18291__A _18263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24229__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23336_ _23336_/CLK _23336_/D VGND VGND VPWR VPWR _13283_/B sky130_fd_sc_hd__dfxtp_4
X_20548_ _20419_/X _20547_/X _24614_/Q _20465_/X VGND VGND VPWR VPWR _20548_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21492__A2 _21638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23267_ _23242_/CLK _23267_/D VGND VGND VPWR VPWR _19631_/A sky130_fd_sc_hd__dfxtp_4
X_20479_ _20461_/X _20478_/Y _15371_/A _20466_/X VGND VGND VPWR VPWR _23708_/D sky130_fd_sc_hd__a2bb2o_4
X_13020_ _13075_/A VGND VGND VPWR VPWR _13299_/A sky130_fd_sc_hd__buf_2
XFILLER_69_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25006_ _25009_/CLK _25006_/D HRESETn VGND VGND VPWR VPWR _25006_/Q sky130_fd_sc_hd__dfrtp_4
X_22218_ _16042_/A _22024_/B _22218_/C _22510_/C VGND VGND VPWR VPWR _22219_/A sky130_fd_sc_hd__or4_4
XFILLER_121_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23198_ _23156_/CLK _19816_/X VGND VGND VPWR VPWR _19812_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_105_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22149_ _24263_/Q _22227_/B VGND VGND VPWR VPWR _22149_/X sky130_fd_sc_hd__and2_4
XFILLER_0_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22526__A1_N _21040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21157__A _17629_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14971_ _14969_/Y _24261_/Q _15224_/A _24258_/Q VGND VGND VPWR VPWR _14971_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23864__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12779__A _22900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16710_ _16710_/A VGND VGND VPWR VPWR _16710_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25088__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13922_ _20710_/B VGND VGND VPWR VPWR _13923_/B sky130_fd_sc_hd__inv_2
X_17690_ _14571_/X _23454_/Q VGND VGND VPWR VPWR _17690_/X sky130_fd_sc_hd__or2_4
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25017__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16641_ _14779_/Y _16639_/X HWDATA[20] _16639_/X VGND VGND VPWR VPWR _16641_/X sky130_fd_sc_hd__a2bb2o_4
X_13853_ _13852_/X VGND VGND VPWR VPWR _14361_/B sky130_fd_sc_hd__inv_2
XFILLER_47_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15631__B1 _15279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12804_ _22778_/A _22779_/A _12802_/Y _12803_/Y VGND VGND VPWR VPWR _12808_/C sky130_fd_sc_hd__o22a_4
X_19360_ _11630_/A VGND VGND VPWR VPWR _19360_/X sky130_fd_sc_hd__buf_2
X_16572_ _14814_/Y _16570_/X _16243_/X _16570_/X VGND VGND VPWR VPWR _24154_/D sky130_fd_sc_hd__a2bb2o_4
X_13784_ _24649_/Q _13761_/A VGND VGND VPWR VPWR _13785_/B sky130_fd_sc_hd__or2_4
XFILLER_43_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18311_ _18290_/X _18311_/B _18310_/Y VGND VGND VPWR VPWR _23855_/D sky130_fd_sc_hd__and3_4
XANTENNA__12996__A1 _12972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15523_ _15503_/X _15504_/X _15522_/X _24548_/Q _15466_/A VGND VGND VPWR VPWR _15523_/X
+ sky130_fd_sc_hd__a32o_4
X_12735_ _12651_/D _12638_/Y VGND VGND VPWR VPWR _12735_/X sky130_fd_sc_hd__or2_4
X_19291_ _23387_/Q VGND VGND VPWR VPWR _21632_/B sky130_fd_sc_hd__inv_2
XFILLER_37_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18242_ _18242_/A _18242_/B _18198_/Y _18257_/B VGND VGND VPWR VPWR _18243_/A sky130_fd_sc_hd__or4_4
X_12666_ _13007_/B VGND VGND VPWR VPWR _12666_/X sky130_fd_sc_hd__buf_2
X_15454_ _15449_/A _15452_/Y _15453_/Y VGND VGND VPWR VPWR _15454_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_8_214_0_HCLK clkbuf_8_215_0_HCLK/A VGND VGND VPWR VPWR _23840_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ _11614_/Y _11610_/X _11616_/X _11610_/X VGND VGND VPWR VPWR _11617_/X sky130_fd_sc_hd__a2bb2o_4
X_14405_ _14383_/A _14383_/B VGND VGND VPWR VPWR _14405_/Y sky130_fd_sc_hd__nand2_4
XFILLER_30_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18173_ _22401_/A _23858_/Q _22401_/A _23858_/Q VGND VGND VPWR VPWR _18177_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24652__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _12650_/A _12595_/Y _12593_/A _12596_/Y VGND VGND VPWR VPWR _12597_/X sky130_fd_sc_hd__a2bb2o_4
X_15385_ _15385_/A VGND VGND VPWR VPWR _22008_/A sky130_fd_sc_hd__inv_2
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17124_ _17053_/A _17124_/B VGND VGND VPWR VPWR _17124_/X sky130_fd_sc_hd__or2_4
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11548_ HWDATA[25] VGND VGND VPWR VPWR _11548_/X sky130_fd_sc_hd__buf_2
X_14336_ _24777_/Q _14325_/X _21549_/A _14327_/X VGND VGND VPWR VPWR _14336_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22680__A1 _24565_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14267_ _13619_/X _18633_/A VGND VGND VPWR VPWR _14273_/A sky130_fd_sc_hd__nor2_4
X_17055_ _17055_/A _17055_/B VGND VGND VPWR VPWR _17055_/X sky130_fd_sc_hd__or2_4
XFILLER_13_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21105__A1_N _17614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24871__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13218_ _13102_/X _13218_/B _13218_/C VGND VGND VPWR VPWR _13218_/X sky130_fd_sc_hd__and3_4
X_16006_ _16014_/A _16014_/B _24359_/Q VGND VGND VPWR VPWR _16006_/X sky130_fd_sc_hd__and3_4
XANTENNA__22432__A1 _24409_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14198_ _20164_/A _20158_/A VGND VGND VPWR VPWR _14198_/X sky130_fd_sc_hd__or2_4
XFILLER_98_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16557__A2_N _16493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13149_ _13110_/A _23324_/Q VGND VGND VPWR VPWR _13150_/C sky130_fd_sc_hd__or2_4
XFILLER_48_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17957_ _17782_/A _17957_/B VGND VGND VPWR VPWR _17957_/X sky130_fd_sc_hd__or2_4
XFILLER_61_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13476__A2 _13480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11593__A HWDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16908_ _16890_/A _16898_/B _16907_/X VGND VGND VPWR VPWR _24074_/D sky130_fd_sc_hd__and3_4
XFILLER_113_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17888_ _17821_/A _17888_/B VGND VGND VPWR VPWR _17888_/X sky130_fd_sc_hd__or2_4
XFILLER_61_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19627_ _21912_/B _19624_/X _19600_/X _19624_/X VGND VGND VPWR VPWR _23269_/D sky130_fd_sc_hd__a2bb2o_4
X_16839_ _16916_/A _16839_/B _16838_/X VGND VGND VPWR VPWR _16840_/B sky130_fd_sc_hd__or3_4
XFILLER_19_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15622__B1 _13658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19558_ _21934_/B _19555_/X _11839_/X _19555_/X VGND VGND VPWR VPWR _23293_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22499__A1 _21870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_24_0_HCLK clkbuf_6_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_49_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18509_ _18509_/A _18509_/B VGND VGND VPWR VPWR _18511_/B sky130_fd_sc_hd__or2_4
XFILLER_0_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19489_ _19488_/Y VGND VGND VPWR VPWR _19489_/X sky130_fd_sc_hd__buf_2
XFILLER_62_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21520_ _21515_/X _21519_/X _21231_/X VGND VGND VPWR VPWR _21528_/B sky130_fd_sc_hd__o21a_4
XFILLER_72_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22626__A _22625_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21451_ _24015_/Q _15653_/X _21448_/X _21449_/X _21450_/X VGND VGND VPWR VPWR _21452_/A
+ sky130_fd_sc_hd__a2111o_4
XANTENNA__24393__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16624__A _16624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20402_ _20402_/A _20212_/B VGND VGND VPWR VPWR _20404_/B sky130_fd_sc_hd__or2_4
XANTENNA__24322__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24170_ _24168_/CLK _16526_/X HRESETn VGND VGND VPWR VPWR _24170_/Q sky130_fd_sc_hd__dfrtp_4
X_21382_ _21385_/A _21382_/B VGND VGND VPWR VPWR _21384_/B sky130_fd_sc_hd__or2_4
XFILLER_135_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22671__B2 _22549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23121_ _23112_/CLK _23121_/D VGND VGND VPWR VPWR _23121_/Q sky130_fd_sc_hd__dfxtp_4
X_20333_ _20249_/A _20333_/B _20332_/Y VGND VGND VPWR VPWR _20333_/X sky130_fd_sc_hd__and3_4
X_23052_ _23036_/X VGND VGND VPWR VPWR IRQ[0] sky130_fd_sc_hd__buf_2
X_20264_ _20264_/A _20264_/B VGND VGND VPWR VPWR _20264_/X sky130_fd_sc_hd__and2_4
XFILLER_103_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22003_ _22306_/A _21976_/X _21983_/X _21997_/X _22002_/X VGND VGND VPWR VPWR _22004_/D
+ sky130_fd_sc_hd__o41a_4
XFILLER_103_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20195_ _20195_/A _20179_/C _20192_/X VGND VGND VPWR VPWR _20195_/X sky130_fd_sc_hd__and3_4
XFILLER_69_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15861__B1 _15772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25181__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19052__B1 _18938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_106_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_213_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12675__B1 _12674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23954_ _23972_/CLK _17584_/Y HRESETn VGND VGND VPWR VPWR _22376_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25110__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21705__A _21793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22905_ _22201_/A _22890_/X _22893_/X _22899_/X _22904_/X VGND VGND VPWR VPWR _22905_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_29_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23885_ _23885_/CLK _18114_/X HRESETn VGND VGND VPWR VPWR _23885_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15613__B1 _24518_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22836_ _22335_/A _22834_/X _22835_/X _24421_/Q _22576_/A VGND VGND VPWR VPWR _22837_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_25_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15422__B _16475_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22767_ _21030_/X _22766_/X _22646_/X _15849_/A _22647_/X VGND VGND VPWR VPWR _22767_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_129_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _12407_/B _12511_/D VGND VGND VPWR VPWR _12520_/Y sky130_fd_sc_hd__nand2_4
X_21718_ _22017_/A VGND VGND VPWR VPWR _22547_/A sky130_fd_sc_hd__buf_2
XFILLER_12_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24506_ _25009_/CLK _24506_/D HRESETn VGND VGND VPWR VPWR _15630_/A sky130_fd_sc_hd__dfrtp_4
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22698_ _22698_/A VGND VGND VPWR VPWR _22698_/Y sky130_fd_sc_hd__inv_2
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _12451_/A _12451_/B VGND VGND VPWR VPWR _12451_/X sky130_fd_sc_hd__or2_4
X_21649_ _22043_/A _21649_/B _21649_/C _20062_/A VGND VGND VPWR VPWR _21649_/X sky130_fd_sc_hd__or4_4
XFILLER_40_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24437_ _24502_/CLK _24437_/D HRESETn VGND VGND VPWR VPWR _22161_/A sky130_fd_sc_hd__dfrtp_4
X_15170_ _15106_/A _15177_/A _15179_/A _15183_/B VGND VGND VPWR VPWR _15170_/X sky130_fd_sc_hd__or4_4
XANTENNA__24063__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12382_ _12382_/A VGND VGND VPWR VPWR _12382_/Y sky130_fd_sc_hd__inv_2
X_24368_ _24425_/CLK _24368_/D HRESETn VGND VGND VPWR VPWR _15981_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22662__B2 _22537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_44_0_HCLK clkbuf_8_45_0_HCLK/A VGND VGND VPWR VPWR _23537_/CLK sky130_fd_sc_hd__clkbuf_1
X_14121_ _14106_/B _14116_/X _14121_/C VGND VGND VPWR VPWR _24850_/D sky130_fd_sc_hd__and3_4
X_23319_ _24750_/CLK _23319_/D VGND VGND VPWR VPWR _23319_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_4_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24299_ _24319_/CLK _24299_/D HRESETn VGND VGND VPWR VPWR _16193_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14052_ _24869_/Q VGND VGND VPWR VPWR _14052_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14989__A _24711_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13003_ _12818_/Y _12999_/X VGND VGND VPWR VPWR _13003_/Y sky130_fd_sc_hd__nand2_4
X_18860_ _18858_/Y _18854_/X _18744_/X _18859_/X VGND VGND VPWR VPWR _18860_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17811_ _17727_/A VGND VGND VPWR VPWR _17944_/A sky130_fd_sc_hd__buf_2
X_18791_ _18789_/Y _18785_/X _18744_/X _18790_/X VGND VGND VPWR VPWR _18791_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15852__B1 _15765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17742_ _17742_/A VGND VGND VPWR VPWR _17899_/A sky130_fd_sc_hd__buf_2
XANTENNA__19043__B1 _19041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14954_ _15136_/C _14960_/A _24660_/Q _14897_/Y VGND VGND VPWR VPWR _14954_/X sky130_fd_sc_hd__a2bb2o_4
X_13905_ _13905_/A VGND VGND VPWR VPWR _13905_/X sky130_fd_sc_hd__buf_2
X_17673_ _14569_/A _17673_/B _17672_/X VGND VGND VPWR VPWR _17673_/X sky130_fd_sc_hd__and3_4
XFILLER_63_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14885_ _24681_/Q VGND VGND VPWR VPWR _14885_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19412_ _19411_/Y _19409_/X _19366_/X _19409_/X VGND VGND VPWR VPWR _19412_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16624_ _16624_/A VGND VGND VPWR VPWR _16624_/X sky130_fd_sc_hd__buf_2
XFILLER_47_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13836_ _13828_/D _13835_/X VGND VGND VPWR VPWR _13880_/C sky130_fd_sc_hd__or2_4
XFILLER_35_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19343_ _13273_/B VGND VGND VPWR VPWR _19343_/Y sky130_fd_sc_hd__inv_2
X_16555_ _16555_/A VGND VGND VPWR VPWR _16555_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24833__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13767_ _13767_/A VGND VGND VPWR VPWR _13797_/A sky130_fd_sc_hd__inv_2
XANTENNA__17250__D _17249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15506_ _15503_/X _15504_/X _15505_/X _24557_/Q _15495_/X VGND VGND VPWR VPWR _24557_/D
+ sky130_fd_sc_hd__a32o_4
X_12718_ _12716_/A _12714_/X _12717_/Y VGND VGND VPWR VPWR _12718_/X sky130_fd_sc_hd__and3_4
X_19274_ _19260_/X VGND VGND VPWR VPWR _19274_/X sky130_fd_sc_hd__buf_2
X_16486_ _16493_/A VGND VGND VPWR VPWR _16486_/X sky130_fd_sc_hd__buf_2
X_13698_ _21733_/A _13687_/X _24918_/Q _13689_/X VGND VGND VPWR VPWR _13698_/X sky130_fd_sc_hd__o22a_4
X_18225_ _23876_/Q _18225_/B VGND VGND VPWR VPWR _18225_/Y sky130_fd_sc_hd__nand2_4
X_15437_ _15436_/Y _14433_/X VGND VGND VPWR VPWR _15437_/X sky130_fd_sc_hd__and2_4
X_12649_ _12629_/X _12584_/Y _12649_/C _12648_/Y VGND VGND VPWR VPWR _12652_/B sky130_fd_sc_hd__or4_4
XANTENNA__12972__A _12972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22165__B _22953_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18156_ _24353_/Q _18234_/A _16050_/Y _18222_/B VGND VGND VPWR VPWR _18163_/A sky130_fd_sc_hd__o22a_4
XANTENNA__18857__B1 _18740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15368_ _11532_/X VGND VGND VPWR VPWR _15368_/X sky130_fd_sc_hd__buf_2
X_17107_ _17042_/D _17096_/B VGND VGND VPWR VPWR _17108_/B sky130_fd_sc_hd__or2_4
XFILLER_50_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11588__A _11599_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14319_ _14315_/C VGND VGND VPWR VPWR _14319_/X sky130_fd_sc_hd__buf_2
XFILLER_32_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18087_ _13050_/A _18085_/X _18086_/Y VGND VGND VPWR VPWR _18087_/X sky130_fd_sc_hd__o21a_4
X_15299_ _15298_/X VGND VGND VPWR VPWR _23762_/D sky130_fd_sc_hd__buf_2
X_17038_ _24042_/Q VGND VGND VPWR VPWR _17040_/A sky130_fd_sc_hd__inv_2
XFILLER_89_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15686__A3 _15494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22405__A1 _11691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22405__B2 _20918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23786__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22612__C _22612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23715__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18989_ _14544_/A _14543_/X _14539_/Y _19904_/D VGND VGND VPWR VPWR _18990_/A sky130_fd_sc_hd__or4_4
XANTENNA__15843__B1 _11545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13308__A _13182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21525__A _21393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20951_ _22087_/A _19550_/Y VGND VGND VPWR VPWR _20953_/B sky130_fd_sc_hd__or2_4
XANTENNA__12133__A2_N _24558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23670_ _23680_/CLK _23670_/D HRESETn VGND VGND VPWR VPWR _17174_/A sky130_fd_sc_hd__dfrtp_4
X_20882_ _20872_/X _20880_/Y _20881_/Y _13381_/Y _11527_/Y VGND VGND VPWR VPWR _20882_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_81_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22621_ _16075_/A _22350_/X _22581_/X VGND VGND VPWR VPWR _22621_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24574__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24503__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22552_ _16343_/Y _21896_/X _16080_/Y _22549_/X VGND VGND VPWR VPWR _22552_/X sky130_fd_sc_hd__o22a_4
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22892__B2 _21187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22356__A _23922_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21503_ _21372_/A _21503_/B _21503_/C VGND VGND VPWR VPWR _21503_/X sky130_fd_sc_hd__and3_4
X_22483_ _22483_/A _20911_/X VGND VGND VPWR VPWR _22483_/X sky130_fd_sc_hd__and2_4
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24222_ _24222_/CLK _24222_/D HRESETn VGND VGND VPWR VPWR _24222_/Q sky130_fd_sc_hd__dfrtp_4
X_21434_ _21434_/A _21430_/X _21433_/X VGND VGND VPWR VPWR _21434_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_3_0_HCLK clkbuf_7_1_0_HCLK/X VGND VGND VPWR VPWR _23246_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_108_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24153_ _24104_/CLK _16574_/X HRESETn VGND VGND VPWR VPWR _24153_/Q sky130_fd_sc_hd__dfrtp_4
X_21365_ _21364_/X VGND VGND VPWR VPWR _21365_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23104_ _23925_/CLK _20068_/X VGND VGND VPWR VPWR _23104_/Q sky130_fd_sc_hd__dfxtp_4
X_20316_ _14257_/Y _20296_/X _20286_/X _20315_/X VGND VGND VPWR VPWR _20317_/A sky130_fd_sc_hd__a211o_4
X_24084_ _24064_/CLK _16873_/X HRESETn VGND VGND VPWR VPWR _24084_/Q sky130_fd_sc_hd__dfrtp_4
X_21296_ _22167_/A _21296_/B _21296_/C VGND VGND VPWR VPWR _21296_/X sky130_fd_sc_hd__and3_4
XFILLER_116_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23035_ _24944_/Q _21703_/B _23033_/X _23034_/Y VGND VGND VPWR VPWR _23035_/X sky130_fd_sc_hd__a211o_4
X_20247_ _20245_/X _20246_/X _15250_/A VGND VGND VPWR VPWR _20247_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21419__B _22155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20178_ _20178_/A VGND VGND VPWR VPWR _20249_/B sky130_fd_sc_hd__inv_2
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13218__A _13102_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21907__B1 _21890_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24986_ _24788_/CLK _13364_/X HRESETn VGND VGND VPWR VPWR _24986_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12112__A2 _24554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21435__A _24096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11951_ _24622_/Q _11951_/B _11512_/Y VGND VGND VPWR VPWR _22510_/B sky130_fd_sc_hd__or3_4
XFILLER_85_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23937_ _23486_/CLK _17659_/X HRESETn VGND VGND VPWR VPWR _13407_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_45_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11961__A _13333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15433__A _16302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11882_ _23785_/Q _11882_/B VGND VGND VPWR VPWR _11894_/A sky130_fd_sc_hd__and2_4
X_14670_ _14625_/A _14625_/B _14625_/A _14625_/B VGND VGND VPWR VPWR _14671_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23868_ _23859_/CLK _23868_/D HRESETn VGND VGND VPWR VPWR _18256_/A sky130_fd_sc_hd__dfrtp_4
X_13621_ _13608_/X _13620_/Y _13330_/X _13620_/Y VGND VGND VPWR VPWR _13621_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15601__A3 _15600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22819_ _22597_/A _22818_/X VGND VGND VPWR VPWR _22819_/X sky130_fd_sc_hd__and2_4
XANTENNA__22332__B1 _22317_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18744__A _18743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23799_ _23796_/CLK _23799_/D HRESETn VGND VGND VPWR VPWR _12039_/A sky130_fd_sc_hd__dfrtp_4
X_16340_ _16338_/Y _16333_/X _16261_/X _16339_/X VGND VGND VPWR VPWR _24241_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24244__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13552_ _13567_/B VGND VGND VPWR VPWR _13580_/A sky130_fd_sc_hd__inv_2
XFILLER_125_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12820__B1 _12818_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12503_ _12379_/Y _12502_/X VGND VGND VPWR VPWR _12503_/X sky130_fd_sc_hd__or2_4
XFILLER_73_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13483_ _13475_/Y _13480_/X _13481_/X _13403_/A _13482_/Y VGND VGND VPWR VPWR _13483_/X
+ sky130_fd_sc_hd__a32o_4
X_16271_ _16268_/X _16269_/X _15494_/X _24271_/Q _16270_/X VGND VGND VPWR VPWR _16271_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16264__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18010_ _17999_/X _15915_/X _18000_/X _23908_/Q _18007_/A VGND VGND VPWR VPWR _23908_/D
+ sky130_fd_sc_hd__a32o_4
X_12434_ _12434_/A _12434_/B _12434_/C VGND VGND VPWR VPWR _25099_/D sky130_fd_sc_hd__and3_4
X_15222_ _15112_/C _15229_/A VGND VGND VPWR VPWR _15222_/X sky130_fd_sc_hd__or2_4
XFILLER_5_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12365_ _12365_/A _12365_/B _12361_/X _12364_/X VGND VGND VPWR VPWR _12365_/X sky130_fd_sc_hd__or4_4
X_15153_ _24673_/Q _15156_/B VGND VGND VPWR VPWR _15153_/X sky130_fd_sc_hd__or2_4
X_14104_ _14104_/A VGND VGND VPWR VPWR _14104_/Y sky130_fd_sc_hd__inv_2
X_15084_ _15083_/X VGND VGND VPWR VPWR _24686_/D sky130_fd_sc_hd__inv_2
X_19961_ _19959_/Y _19960_/X _19387_/X _19960_/X VGND VGND VPWR VPWR _19961_/X sky130_fd_sc_hd__a2bb2o_4
X_12296_ _12265_/B _12300_/A VGND VGND VPWR VPWR _12297_/B sky130_fd_sc_hd__nand2_4
XFILLER_5_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12841__A1_N _12947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14035_ _20221_/B _14026_/X _13632_/X _14028_/X VGND VGND VPWR VPWR _14035_/X sky130_fd_sc_hd__a2bb2o_4
X_18912_ _23521_/Q VGND VGND VPWR VPWR _18912_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19892_ _23171_/Q VGND VGND VPWR VPWR _21673_/B sky130_fd_sc_hd__inv_2
XANTENNA__19264__B1 _19149_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21071__B1 _20782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25032__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18843_ _21506_/B _18838_/X _15559_/X _18838_/X VGND VGND VPWR VPWR _18843_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18919__A _17684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18774_ _18773_/Y _18769_/X _18679_/X _18769_/X VGND VGND VPWR VPWR _23570_/D sky130_fd_sc_hd__a2bb2o_4
X_15986_ _24366_/Q VGND VGND VPWR VPWR _15986_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17725_ _17725_/A VGND VGND VPWR VPWR _17738_/A sky130_fd_sc_hd__buf_2
X_14937_ _24260_/Q VGND VGND VPWR VPWR _14937_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17656_ _15810_/B _17655_/X VGND VGND VPWR VPWR _17656_/Y sky130_fd_sc_hd__nor2_4
X_14868_ _14702_/Y _14868_/B VGND VGND VPWR VPWR _14879_/C sky130_fd_sc_hd__or2_4
XANTENNA__16250__B1 _24280_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16607_ _14816_/Y _16606_/X _16455_/X _16606_/X VGND VGND VPWR VPWR _24133_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13819_ _13828_/A _13867_/A _13867_/C VGND VGND VPWR VPWR _13851_/B sky130_fd_sc_hd__or3_4
X_17587_ _17484_/Y _17587_/B VGND VGND VPWR VPWR _17587_/X sky130_fd_sc_hd__or2_4
XFILLER_56_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14799_ _15045_/A _16594_/A _15045_/A _16594_/A VGND VGND VPWR VPWR _14799_/X sky130_fd_sc_hd__a2bb2o_4
X_19326_ _19799_/A _18064_/X _18666_/C VGND VGND VPWR VPWR _19327_/A sky130_fd_sc_hd__or3_4
XFILLER_17_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16538_ _16537_/Y _16535_/X _16369_/X _16535_/X VGND VGND VPWR VPWR _16538_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16002__B1 _15291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19257_ _20978_/B _19251_/X _19256_/X _19238_/Y VGND VGND VPWR VPWR _19257_/X sky130_fd_sc_hd__a2bb2o_4
X_16469_ _24192_/Q VGND VGND VPWR VPWR _16469_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16174__A _24306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18208_ _23858_/Q VGND VGND VPWR VPWR _18295_/A sky130_fd_sc_hd__inv_2
X_19188_ _23422_/Q VGND VGND VPWR VPWR _19188_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23967__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18139_ _23855_/Q VGND VGND VPWR VPWR _18213_/D sky130_fd_sc_hd__inv_2
XFILLER_89_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22623__B _22435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21150_ _21130_/A VGND VGND VPWR VPWR _21155_/A sky130_fd_sc_hd__buf_2
XFILLER_137_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_90_0_HCLK clkbuf_8_91_0_HCLK/A VGND VGND VPWR VPWR _23618_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16621__B _16235_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20101_ _21931_/B _20098_/X _19600_/A _20098_/X VGND VGND VPWR VPWR _20101_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22929__A2 _22311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21081_ _21113_/B VGND VGND VPWR VPWR _21082_/B sky130_fd_sc_hd__buf_2
XFILLER_63_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16069__B1 _15765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20032_ _20947_/B _20027_/X _19755_/X _20014_/Y VGND VGND VPWR VPWR _20032_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11765__B _11728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17733__A _17727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24840_ _24840_/CLK _24840_/D HRESETn VGND VGND VPWR VPWR _23042_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21551__A1_N _14255_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12072__A2_N _24556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19558__B2 _19555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21983_ _21978_/X _21982_/X VGND VGND VPWR VPWR _21983_/X sky130_fd_sc_hd__and2_4
XFILLER_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24755__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24771_ _24897_/CLK _24771_/D HRESETn VGND VGND VPWR VPWR scl_oen_o_S4 sky130_fd_sc_hd__dfstp_4
XFILLER_6_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11781__A _11694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20934_ _20931_/X _20933_/X _24964_/Q _22439_/B VGND VGND VPWR VPWR _20935_/A sky130_fd_sc_hd__o22a_4
X_23722_ _23744_/CLK _23722_/D HRESETn VGND VGND VPWR VPWR _20534_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20865_ _20806_/A VGND VGND VPWR VPWR _20866_/A sky130_fd_sc_hd__buf_2
XPHY_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23653_ _23852_/CLK _23653_/D HRESETn VGND VGND VPWR VPWR _20735_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__15595__A2 _15582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22604_ _21040_/X _22600_/Y _22601_/X _22603_/X VGND VGND VPWR VPWR _22604_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23584_ _23586_/CLK _18729_/X VGND VGND VPWR VPWR _17920_/B sky130_fd_sc_hd__dfxtp_4
X_20796_ _20806_/A VGND VGND VPWR VPWR _21285_/B sky130_fd_sc_hd__buf_2
XPHY_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22535_ _22500_/Y _22509_/X _22661_/C _22534_/X VGND VGND VPWR VPWR HRDATA[16] sky130_fd_sc_hd__or4_4
XFILLER_127_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14555__B1 _13462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22617__A1 _24274_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22466_ _16181_/A _22246_/B VGND VGND VPWR VPWR _22466_/X sky130_fd_sc_hd__or2_4
XFILLER_10_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21417_ _21410_/X _21416_/X _21062_/X VGND VGND VPWR VPWR _21538_/A sky130_fd_sc_hd__o21a_4
X_24205_ _24244_/CLK _16437_/X HRESETn VGND VGND VPWR VPWR _24205_/Q sky130_fd_sc_hd__dfrtp_4
X_25185_ _24847_/CLK _25185_/D HRESETn VGND VGND VPWR VPWR _25185_/Q sky130_fd_sc_hd__dfrtp_4
X_22397_ _12498_/A _22178_/X _24040_/Q _22260_/X VGND VGND VPWR VPWR _22398_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12117__A _12117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23637__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16812__A _17132_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12150_ _25124_/Q _12148_/Y _12149_/Y _24565_/Q VGND VGND VPWR VPWR _12150_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14307__B1 _14218_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24136_ _24145_/CLK _16603_/X HRESETn VGND VGND VPWR VPWR _16601_/A sky130_fd_sc_hd__dfrtp_4
X_21348_ _21348_/A _19700_/Y VGND VGND VPWR VPWR _21350_/B sky130_fd_sc_hd__or2_4
Xclkbuf_8_118_0_HCLK clkbuf_7_59_0_HCLK/X VGND VGND VPWR VPWR _24644_/CLK sky130_fd_sc_hd__clkbuf_1
X_12081_ _12081_/A _12081_/B _12077_/X _12081_/D VGND VGND VPWR VPWR _12120_/A sky130_fd_sc_hd__or4_4
XANTENNA__15428__A _21179_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24067_ _24620_/CLK _16936_/X HRESETn VGND VGND VPWR VPWR _24067_/Q sky130_fd_sc_hd__dfrtp_4
X_21279_ _23023_/A _21274_/X _21279_/C VGND VGND VPWR VPWR _21324_/A sky130_fd_sc_hd__and3_4
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23067__D _20550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23018_ _24156_/Q _22505_/A _22840_/X _23017_/X VGND VGND VPWR VPWR _23019_/C sky130_fd_sc_hd__a211o_4
XFILLER_81_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18739__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15840_ _15839_/Y _15834_/X _15756_/X _15834_/X VGND VGND VPWR VPWR _24422_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23626__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19549__B2 _19546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21165__A _21153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15771_ _12851_/Y _15768_/X _15770_/X _15768_/X VGND VGND VPWR VPWR _24449_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24496__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12983_ _12805_/Y _12992_/B VGND VGND VPWR VPWR _12984_/B sky130_fd_sc_hd__or2_4
X_24969_ _24750_/CLK _24969_/D HRESETn VGND VGND VPWR VPWR _13468_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16259__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17510_ _16746_/X _17510_/B VGND VGND VPWR VPWR _17511_/B sky130_fd_sc_hd__and2_4
X_14722_ _14722_/A VGND VGND VPWR VPWR _14722_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11934_ _11933_/Y _11931_/X _20880_/A _11931_/X VGND VGND VPWR VPWR _11934_/X sky130_fd_sc_hd__a2bb2o_4
X_18490_ _23834_/Q _18489_/Y VGND VGND VPWR VPWR _18492_/B sky130_fd_sc_hd__or2_4
XANTENNA__24425__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17441_ _17408_/D VGND VGND VPWR VPWR _17441_/Y sky130_fd_sc_hd__inv_2
X_14653_ _24725_/Q _14612_/X _24725_/Q _14612_/X VGND VGND VPWR VPWR _14653_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11865_ _11649_/Y _13551_/B _11708_/A _11645_/X VGND VGND VPWR VPWR _11871_/D sky130_fd_sc_hd__a211o_4
XANTENNA__15586__A2 _15582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13604_ _11676_/A _11683_/A VGND VGND VPWR VPWR _13604_/X sky130_fd_sc_hd__or2_4
X_17372_ _17313_/X _17371_/X VGND VGND VPWR VPWR _17373_/B sky130_fd_sc_hd__or2_4
X_11796_ _11803_/C _11796_/B VGND VGND VPWR VPWR _11796_/Y sky130_fd_sc_hd__nor2_4
X_14584_ _24733_/Q VGND VGND VPWR VPWR _14596_/A sky130_fd_sc_hd__inv_2
XFILLER_41_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19111_ _17845_/B VGND VGND VPWR VPWR _19111_/Y sky130_fd_sc_hd__inv_2
X_16323_ _24247_/Q VGND VGND VPWR VPWR _16323_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20867__B1 _24093_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13535_ _23738_/Q _20599_/A _13535_/C _20611_/A VGND VGND VPWR VPWR _13535_/X sky130_fd_sc_hd__or4_4
XANTENNA__14507__A _14506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19042_ _19034_/Y VGND VGND VPWR VPWR _19042_/X sky130_fd_sc_hd__buf_2
X_16254_ HWDATA[22] VGND VGND VPWR VPWR _16254_/X sky130_fd_sc_hd__buf_2
XFILLER_71_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13466_ _13463_/Y VGND VGND VPWR VPWR _13480_/A sky130_fd_sc_hd__buf_2
XFILLER_16_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15205_ _14883_/Y _15207_/B _15204_/Y VGND VGND VPWR VPWR _24661_/D sky130_fd_sc_hd__o21a_4
XFILLER_51_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12417_ _12417_/A _12417_/B VGND VGND VPWR VPWR _12424_/A sky130_fd_sc_hd__or2_4
XFILLER_138_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16185_ _16183_/Y _16178_/X _15369_/X _16184_/X VGND VGND VPWR VPWR _24303_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19485__B1 _19392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13397_ _16302_/A _13328_/X VGND VGND VPWR VPWR _13397_/Y sky130_fd_sc_hd__nor2_4
XFILLER_12_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23010__A1_N _21546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16722__A _23947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_14_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__25213__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15136_ _15159_/A _15159_/B _15136_/C _15115_/A VGND VGND VPWR VPWR _15152_/A sky130_fd_sc_hd__or4_4
X_12348_ _12348_/A VGND VGND VPWR VPWR _12534_/A sky130_fd_sc_hd__inv_2
XFILLER_86_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_77_0_HCLK clkbuf_7_76_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_77_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12279_ _12097_/Y _12282_/B VGND VGND VPWR VPWR _12279_/Y sky130_fd_sc_hd__nand2_4
X_15067_ _14743_/X _15067_/B _15067_/C _15079_/B VGND VGND VPWR VPWR _15067_/X sky130_fd_sc_hd__or4_4
X_19944_ _19943_/Y _19939_/X _19859_/X _19926_/Y VGND VGND VPWR VPWR _23151_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23033__B2 _20919_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14018_ _11951_/B VGND VGND VPWR VPWR _15314_/B sky130_fd_sc_hd__inv_2
XANTENNA__16466__A1_N _16464_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19875_ _19875_/A VGND VGND VPWR VPWR _21392_/B sky130_fd_sc_hd__inv_2
XFILLER_68_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22792__B1 _14913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17553__A _16692_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18826_ _18825_/Y _18822_/X _18802_/X _18822_/X VGND VGND VPWR VPWR _18826_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18757_ _18756_/Y _18752_/X _18712_/X _18752_/A VGND VGND VPWR VPWR _18757_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15969_ _15968_/Y _15966_/X _11590_/X _15966_/X VGND VGND VPWR VPWR _15969_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22544__B1 _14751_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16169__A _24308_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17708_ _17705_/X VGND VGND VPWR VPWR _17708_/X sky130_fd_sc_hd__buf_2
XANTENNA__24166__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18688_ _18687_/Y _18682_/X _16556_/X _18682_/A VGND VGND VPWR VPWR _18688_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_58_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17639_ _17639_/A VGND VGND VPWR VPWR _17639_/X sky130_fd_sc_hd__buf_2
X_20650_ _20648_/Y _20644_/X _20649_/X VGND VGND VPWR VPWR _20650_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15801__A _15801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20419__A _20511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19309_ _19307_/Y _19305_/X _19308_/X _19305_/X VGND VGND VPWR VPWR _19309_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20858__B1 _22153_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19712__B2 _19710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20581_ _16539_/Y _20574_/X _20562_/X _20580_/Y VGND VGND VPWR VPWR _20582_/A sky130_fd_sc_hd__o22a_4
X_22320_ _20917_/X _22318_/X _20903_/X _22319_/X VGND VGND VPWR VPWR _22320_/X sky130_fd_sc_hd__o22a_4
XFILLER_34_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22634__A _22629_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22251_ _22835_/A VGND VGND VPWR VPWR _22251_/X sky130_fd_sc_hd__buf_2
XFILLER_30_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19476__B1 _19381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23730__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21202_ _21202_/A VGND VGND VPWR VPWR _21372_/A sky130_fd_sc_hd__buf_2
X_22182_ _22182_/A _22181_/X VGND VGND VPWR VPWR _22182_/X sky130_fd_sc_hd__and2_4
X_21133_ _21153_/A VGND VGND VPWR VPWR _21352_/A sky130_fd_sc_hd__buf_2
XANTENNA__19228__B1 _19227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23024__B2 _22531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21064_ _15821_/X VGND VGND VPWR VPWR _21064_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24936__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11523__B1 _11522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20015_ _20014_/Y VGND VGND VPWR VPWR _20015_/X sky130_fd_sc_hd__buf_2
XFILLER_8_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_28_0_HCLK_A clkbuf_4_14_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15804__A3 _15735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24823_ _24823_/CLK _14203_/X HRESETn VGND VGND VPWR VPWR _20195_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21889__A2 _13335_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19400__B1 _19308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24754_ _24757_/CLK _24754_/D HRESETn VGND VGND VPWR VPWR _14424_/A sky130_fd_sc_hd__dfrtp_4
X_21966_ _14494_/X _21945_/Y _21952_/Y _21959_/Y _21965_/Y VGND VGND VPWR VPWR _21967_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_54_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16214__B1 _15801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23705_ _23706_/CLK _20467_/X HRESETn VGND VGND VPWR VPWR _23705_/Q sky130_fd_sc_hd__dfrtp_4
X_20917_ _13609_/X VGND VGND VPWR VPWR _20917_/X sky130_fd_sc_hd__buf_2
XPHY_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ _21897_/A _21106_/X VGND VGND VPWR VPWR _21897_/X sky130_fd_sc_hd__and2_4
XPHY_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24685_ _24681_/CLK _15089_/X HRESETn VGND VGND VPWR VPWR _14785_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11650_/A VGND VGND VPWR VPWR _13557_/A sky130_fd_sc_hd__inv_2
XPHY_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ _17217_/Y _13614_/X _24914_/Q _21093_/B VGND VGND VPWR VPWR _20849_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23636_ _23641_/CLK _23636_/D HRESETn VGND VGND VPWR VPWR _18614_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23889__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11581_ _16087_/A VGND VGND VPWR VPWR _11581_/X sky130_fd_sc_hd__buf_2
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20779_ _22933_/B VGND VGND VPWR VPWR _20780_/A sky130_fd_sc_hd__buf_2
XFILLER_80_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23567_ _23586_/CLK _23567_/D VGND VGND VPWR VPWR _17956_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23818__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13320_ _11710_/X _13304_/X _13319_/X _24997_/Q _11708_/X VGND VGND VPWR VPWR _13320_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22518_ _24445_/Q _21979_/X VGND VGND VPWR VPWR _22518_/X sky130_fd_sc_hd__or2_4
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23498_ _23586_/CLK _23498_/D VGND VGND VPWR VPWR _13197_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13251_ _13219_/A _13251_/B VGND VGND VPWR VPWR _13251_/X sky130_fd_sc_hd__or2_4
X_22449_ _22449_/A _20802_/X VGND VGND VPWR VPWR _22449_/X sky130_fd_sc_hd__and2_4
XFILLER_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16542__A _16530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12202_ _12190_/A _12200_/X _12201_/X VGND VGND VPWR VPWR _25131_/D sky130_fd_sc_hd__and3_4
X_13182_ _13182_/A _19380_/A VGND VGND VPWR VPWR _13182_/X sky130_fd_sc_hd__or2_4
XANTENNA__12594__A2_N _12592_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25168_ _23898_/CLK _25168_/D HRESETn VGND VGND VPWR VPWR _13053_/A sky130_fd_sc_hd__dfrtp_4
X_12133_ _12132_/Y _24558_/Q _12132_/Y _24558_/Q VGND VGND VPWR VPWR _12133_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15158__A _15158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19219__B1 _19152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24119_ _24112_/CLK _24119_/D HRESETn VGND VGND VPWR VPWR _22857_/A sky130_fd_sc_hd__dfrtp_4
X_17990_ _15430_/A VGND VGND VPWR VPWR _17990_/X sky130_fd_sc_hd__buf_2
X_25099_ _23716_/CLK _25099_/D HRESETn VGND VGND VPWR VPWR _12432_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17076__C _17053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12064_ _12063_/X VGND VGND VPWR VPWR _12065_/A sky130_fd_sc_hd__buf_2
X_16941_ _16937_/B _16941_/B _16951_/C VGND VGND VPWR VPWR _16941_/X sky130_fd_sc_hd__and3_4
XFILLER_96_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24677__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21577__B2 _21020_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14997__A _14997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19660_ _19658_/Y _19659_/X _19614_/X _19659_/X VGND VGND VPWR VPWR _23257_/D sky130_fd_sc_hd__a2bb2o_4
X_16872_ _16863_/A _16875_/B _16849_/X VGND VGND VPWR VPWR _16872_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24606__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18611_ _20292_/A _20289_/A VGND VGND VPWR VPWR _20293_/A sky130_fd_sc_hd__or2_4
XANTENNA__16453__B1 _16451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15823_ _15822_/X VGND VGND VPWR VPWR _16135_/B sky130_fd_sc_hd__inv_2
X_19591_ _21223_/B _19588_/X _19462_/X _19588_/X VGND VGND VPWR VPWR _23280_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18542_ _18540_/A _18536_/B _18541_/Y VGND VGND VPWR VPWR _18542_/X sky130_fd_sc_hd__and3_4
X_15754_ _12813_/Y _15752_/X _15753_/X _15752_/X VGND VGND VPWR VPWR _24458_/D sky130_fd_sc_hd__a2bb2o_4
X_12966_ _22396_/A _12965_/Y VGND VGND VPWR VPWR _12966_/X sky130_fd_sc_hd__or2_4
X_14705_ _14696_/X _14698_/X _14705_/C _14704_/X VGND VGND VPWR VPWR _14705_/X sky130_fd_sc_hd__or4_4
X_11917_ _13391_/B _11916_/X _24976_/Q _11917_/D VGND VGND VPWR VPWR _11918_/A sky130_fd_sc_hd__or4_4
X_18473_ _18416_/Y _18470_/X VGND VGND VPWR VPWR _18473_/X sky130_fd_sc_hd__or2_4
X_15685_ _15664_/A VGND VGND VPWR VPWR _15685_/X sky130_fd_sc_hd__buf_2
X_12897_ _12860_/Y _12894_/X _12888_/Y _12896_/X VGND VGND VPWR VPWR _12898_/A sky130_fd_sc_hd__a211o_4
XFILLER_61_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17424_ _17317_/C _17412_/B VGND VGND VPWR VPWR _17425_/C sky130_fd_sc_hd__nand2_4
XANTENNA__15621__A _15604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14636_ _14655_/A VGND VGND VPWR VPWR _14636_/X sky130_fd_sc_hd__buf_2
XFILLER_18_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11848_ _19607_/A VGND VGND VPWR VPWR _11848_/X sky130_fd_sc_hd__buf_2
XANTENNA__22829__B2 _22657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17355_ _17329_/A _17327_/X _17305_/Y VGND VGND VPWR VPWR _17355_/X sky130_fd_sc_hd__o21a_4
X_14567_ _17674_/A VGND VGND VPWR VPWR _17732_/A sky130_fd_sc_hd__buf_2
XFILLER_18_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11779_ _25180_/Q _11828_/B _11769_/A VGND VGND VPWR VPWR _11784_/B sky130_fd_sc_hd__or3_4
XANTENNA__18932__A _18678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16306_ _16305_/X _16306_/B VGND VGND VPWR VPWR _16313_/A sky130_fd_sc_hd__nor2_4
XANTENNA__13141__A _13316_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13518_ _23066_/Q _13517_/Y VGND VGND VPWR VPWR _13518_/X sky130_fd_sc_hd__and2_4
X_17286_ _23998_/Q VGND VGND VPWR VPWR _17286_/Y sky130_fd_sc_hd__inv_2
X_14498_ _21403_/A _14506_/B _14484_/X _14497_/X VGND VGND VPWR VPWR _14498_/X sky130_fd_sc_hd__o22a_4
X_19025_ _19012_/Y VGND VGND VPWR VPWR _19025_/X sky130_fd_sc_hd__buf_2
X_16237_ _16237_/A VGND VGND VPWR VPWR _16237_/X sky130_fd_sc_hd__buf_2
XFILLER_16_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19775__A2_N _19772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13449_ _13449_/A VGND VGND VPWR VPWR _14387_/C sky130_fd_sc_hd__buf_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16168_ _16167_/Y _16165_/X _15770_/X _16165_/X VGND VGND VPWR VPWR _16168_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11596__A _25201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15119_ _15118_/X VGND VGND VPWR VPWR _15119_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23006__A1 _23026_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23006__B2 _22460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16099_ _16084_/A VGND VGND VPWR VPWR _16099_/X sky130_fd_sc_hd__buf_2
XFILLER_114_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19927_ _19926_/Y VGND VGND VPWR VPWR _19927_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_101_0_HCLK clkbuf_7_50_0_HCLK/X VGND VGND VPWR VPWR _24859_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__13401__A1_N _20883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21568__A1 _24549_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_164_0_HCLK clkbuf_7_82_0_HCLK/X VGND VGND VPWR VPWR _23489_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_69_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24347__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_7_0_HCLK clkbuf_7_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19858_ _19858_/A VGND VGND VPWR VPWR _21002_/B sky130_fd_sc_hd__inv_2
XFILLER_68_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14700__A _14997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16444__B1 _16096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18809_ _18809_/A VGND VGND VPWR VPWR _18809_/X sky130_fd_sc_hd__buf_2
XFILLER_3_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19789_ _19788_/Y _19786_/X _19452_/X _19786_/X VGND VGND VPWR VPWR _23211_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13316__A _13316_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21820_ _20967_/A _21818_/X _21820_/C VGND VGND VPWR VPWR _21820_/X sky130_fd_sc_hd__and3_4
XFILLER_37_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22629__A _22629_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21751_ _21751_/A _19276_/Y VGND VGND VPWR VPWR _21752_/C sky130_fd_sc_hd__or2_4
XFILLER_92_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16627__A _16627_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20702_ _20702_/A VGND VGND VPWR VPWR _20703_/B sky130_fd_sc_hd__inv_2
XANTENNA__15531__A _16302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21740__B2 _20866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21682_ _21665_/A _21680_/X _21681_/X VGND VGND VPWR VPWR _21682_/X sky130_fd_sc_hd__and3_4
XANTENNA__21252__B _20827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24470_ _24478_/CLK _15707_/X HRESETn VGND VGND VPWR VPWR _24470_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23982__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12874__B _12818_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20633_ _20621_/X _20632_/Y _24175_/Q _20624_/X VGND VGND VPWR VPWR _23744_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23421_ _23596_/CLK _19194_/X VGND VGND VPWR VPWR _23421_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23911__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25135__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23352_ _23336_/CLK _23352_/D VGND VGND VPWR VPWR _19389_/A sky130_fd_sc_hd__dfxtp_4
X_20564_ _16551_/Y _20553_/X _20562_/X _20563_/X VGND VGND VPWR VPWR _20564_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22364__A _20753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22303_ _24478_/Q _22999_/B VGND VGND VPWR VPWR _22303_/X sky130_fd_sc_hd__or2_4
X_23283_ _23282_/CLK _23283_/D VGND VGND VPWR VPWR _19583_/A sky130_fd_sc_hd__dfxtp_4
X_20495_ _20495_/A _20495_/B _20495_/C VGND VGND VPWR VPWR _20495_/X sky130_fd_sc_hd__and3_4
XANTENNA__22083__B _20918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22234_ _22225_/X _22229_/X _22231_/X _22233_/X VGND VGND VPWR VPWR _22235_/B sky130_fd_sc_hd__o22a_4
XANTENNA__14698__A2_N _24124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25022_ _24566_/CLK _12952_/X HRESETn VGND VGND VPWR VPWR _12951_/A sky130_fd_sc_hd__dfrtp_4
X_22165_ _16198_/A _22953_/B VGND VGND VPWR VPWR _22165_/X sky130_fd_sc_hd__and2_4
XANTENNA__19673__A _19680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_60_0_HCLK clkbuf_7_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_60_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21116_ _13391_/A _20872_/X _11933_/Y _11960_/A VGND VGND VPWR VPWR _21116_/X sky130_fd_sc_hd__o22a_4
XFILLER_120_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22096_ _20962_/A _22094_/X _22095_/X VGND VGND VPWR VPWR _22096_/X sky130_fd_sc_hd__and3_4
X_21047_ _21047_/A VGND VGND VPWR VPWR _21047_/X sky130_fd_sc_hd__buf_2
XANTENNA__15706__A _11630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24088__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22220__A2 _20927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16435__B1 _16179_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24017__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22508__B1 _23023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12820_ _25007_/Q _21269_/A _12818_/Y _12819_/Y VGND VGND VPWR VPWR _12821_/D sky130_fd_sc_hd__o22a_4
X_24806_ _23774_/CLK _14251_/X HRESETn VGND VGND VPWR VPWR _24806_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22998_ _22978_/X _22982_/X _22997_/X VGND VGND VPWR VPWR HRDATA[30] sky130_fd_sc_hd__a21o_4
X_12751_ _12749_/A _12742_/B _12751_/C VGND VGND VPWR VPWR _12751_/X sky130_fd_sc_hd__and3_4
XFILLER_61_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24737_ _24735_/CLK _24737_/D HRESETn VGND VGND VPWR VPWR _14563_/A sky130_fd_sc_hd__dfrtp_4
X_21949_ _21374_/A _21949_/B VGND VGND VPWR VPWR _21951_/B sky130_fd_sc_hd__or2_4
XPHY_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21731__A1 _20819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _11696_/X _11702_/B VGND VGND VPWR VPWR _11702_/X sky130_fd_sc_hd__or2_4
XANTENNA__15441__A _15439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14983__C _14990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15464_/X VGND VGND VPWR VPWR _15470_/Y sky130_fd_sc_hd__inv_2
XPHY_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12547_/Y _12679_/X VGND VGND VPWR VPWR _12683_/C sky130_fd_sc_hd__or2_4
XPHY_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24668_ _24671_/CLK _24668_/D HRESETn VGND VGND VPWR VPWR _24668_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _14419_/Y _14420_/X _14412_/X _14415_/X _14420_/A VGND VGND VPWR VPWR _24756_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_42_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _25192_/Q VGND VGND VPWR VPWR _11633_/Y sky130_fd_sc_hd__inv_2
XPHY_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23619_ _24788_/CLK _20701_/X HRESETn VGND VGND VPWR VPWR _20269_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__23652__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14057__A _24867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24599_ _23706_/CLK _15367_/X HRESETn VGND VGND VPWR VPWR _24599_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17140_ _17034_/C _17134_/X VGND VGND VPWR VPWR _17153_/B sky130_fd_sc_hd__or2_4
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14352_ _14352_/A _14357_/B _14352_/C _13841_/X VGND VGND VPWR VPWR _14353_/A sky130_fd_sc_hd__or4_4
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11564_ _11562_/Y _11559_/X _11563_/X _11559_/X VGND VGND VPWR VPWR _11564_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13303_ _13271_/A _13303_/B _13303_/C VGND VGND VPWR VPWR _13304_/C sky130_fd_sc_hd__or3_4
XFILLER_6_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17071_ _17052_/A _17069_/X _17070_/X VGND VGND VPWR VPWR _17071_/X sky130_fd_sc_hd__and3_4
X_14283_ _14282_/Y _14280_/X _14094_/X _14280_/X VGND VGND VPWR VPWR _24793_/D sky130_fd_sc_hd__a2bb2o_4
X_16022_ _17806_/A VGND VGND VPWR VPWR _16022_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21247__B1 _21246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13234_ _13202_/A _13234_/B VGND VGND VPWR VPWR _13235_/C sky130_fd_sc_hd__or2_4
XANTENNA__24858__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22995__B1 _22407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13165_ _13127_/A _23073_/Q VGND VGND VPWR VPWR _13167_/B sky130_fd_sc_hd__or2_4
XANTENNA__16674__B1 _24093_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12116_ _12116_/A VGND VGND VPWR VPWR _12174_/A sky130_fd_sc_hd__inv_2
X_13096_ _11741_/X VGND VGND VPWR VPWR _13244_/A sky130_fd_sc_hd__buf_2
X_17973_ _16231_/A _11720_/X VGND VGND VPWR VPWR _17973_/X sky130_fd_sc_hd__or2_4
XFILLER_46_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12047_ _20697_/B VGND VGND VPWR VPWR _20695_/B sky130_fd_sc_hd__buf_2
X_16924_ _16831_/D _16924_/B VGND VGND VPWR VPWR _16937_/B sky130_fd_sc_hd__or2_4
X_19712_ _22091_/B _19710_/X _19711_/X _19710_/X VGND VGND VPWR VPWR _23238_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24440__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_237_0_HCLK clkbuf_8_237_0_HCLK/A VGND VGND VPWR VPWR _24177_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16855_ _16774_/A _16854_/Y VGND VGND VPWR VPWR _16855_/X sky130_fd_sc_hd__or2_4
X_19643_ _19643_/A VGND VGND VPWR VPWR _22110_/B sky130_fd_sc_hd__inv_2
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16142__A2_N _16138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18927__A _18935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15806_ _15807_/A _13456_/A VGND VGND VPWR VPWR _15806_/Y sky130_fd_sc_hd__nor2_4
XFILLER_65_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13136__A _13136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19574_ _14544_/A _14543_/X _14493_/X _19904_/D VGND VGND VPWR VPWR _19575_/A sky130_fd_sc_hd__or4_4
XFILLER_92_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16786_ _24060_/Q VGND VGND VPWR VPWR _16921_/C sky130_fd_sc_hd__inv_2
XFILLER_98_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13998_ _13925_/C _13998_/B VGND VGND VPWR VPWR _13999_/A sky130_fd_sc_hd__or2_4
XFILLER_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18525_ _18421_/B _18545_/A VGND VGND VPWR VPWR _18543_/B sky130_fd_sc_hd__or2_4
XFILLER_98_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15737_ _15582_/X _15641_/X _15735_/X _20738_/B _15736_/X VGND VGND VPWR VPWR _15737_/X
+ sky130_fd_sc_hd__a32o_4
X_12949_ _12952_/A _12943_/X _12949_/C VGND VGND VPWR VPWR _12949_/X sky130_fd_sc_hd__and3_4
XANTENNA__16729__B2 _16692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13660__B1 _11604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18456_ _18463_/A _18454_/X _18455_/X VGND VGND VPWR VPWR _23842_/D sky130_fd_sc_hd__and3_4
X_15668_ _12380_/Y _15666_/X _15332_/X _15666_/X VGND VGND VPWR VPWR _24495_/D sky130_fd_sc_hd__a2bb2o_4
X_17407_ _17303_/Y _17323_/D VGND VGND VPWR VPWR _17408_/D sky130_fd_sc_hd__or2_4
X_14619_ _14619_/A VGND VGND VPWR VPWR _14620_/A sky130_fd_sc_hd__buf_2
XFILLER_21_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18387_ _16441_/Y _18517_/A _16441_/Y _18517_/A VGND VGND VPWR VPWR _18387_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15599_ _15740_/A VGND VGND VPWR VPWR _15599_/X sky130_fd_sc_hd__buf_2
XANTENNA__18662__A _19859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17338_ _17338_/A VGND VGND VPWR VPWR _17338_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22184__A _12346_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11974__B1 _11626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17269_ _17269_/A _17269_/B _17259_/X _17269_/D VGND VGND VPWR VPWR _17297_/A sky130_fd_sc_hd__or4_4
X_19008_ _20990_/B _19003_/X _18662_/X _18990_/Y VGND VGND VPWR VPWR _19008_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20280_ _14241_/Y _20273_/X _14266_/X _20279_/X VGND VGND VPWR VPWR _20281_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24599__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24528__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_47_0_HCLK clkbuf_6_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_95_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16665__B1 _16369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16725__A2_N _22434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21528__A _21396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24181__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23970_ _24361_/CLK _17522_/Y HRESETn VGND VGND VPWR VPWR _22920_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_60_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16417__B1 _15484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24110__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22921_ _22921_/A _22418_/X VGND VGND VPWR VPWR _22921_/X sky130_fd_sc_hd__and2_4
XFILLER_42_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17741__A _17732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20544__A1_N _20419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22852_ _22852_/A VGND VGND VPWR VPWR _23004_/A sky130_fd_sc_hd__buf_2
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_21803_ _21802_/X VGND VGND VPWR VPWR _21803_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21263__A _12349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12454__A1 _12448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17460__B _17460_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13651__B1 _11585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22783_ _22783_/A _22505_/A VGND VGND VPWR VPWR _22783_/X sky130_fd_sc_hd__and2_4
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24522_ _24523_/CLK _24522_/D HRESETn VGND VGND VPWR VPWR _24522_/Q sky130_fd_sc_hd__dfrtp_4
X_21734_ _20246_/A _21638_/X _14083_/A _21179_/A VGND VGND VPWR VPWR _21734_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19668__A _19680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24453_ _24432_/CLK _15762_/X HRESETn VGND VGND VPWR VPWR _22779_/A sky130_fd_sc_hd__dfrtp_4
X_21665_ _21665_/A _21663_/X _21664_/X VGND VGND VPWR VPWR _21665_/X sky130_fd_sc_hd__and3_4
XANTENNA__22806__B _22806_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23404_ _23939_/CLK _23404_/D VGND VGND VPWR VPWR _19243_/A sky130_fd_sc_hd__dfxtp_4
X_20616_ _20598_/X _20615_/Y _16522_/A _20603_/X VGND VGND VPWR VPWR _20616_/X sky130_fd_sc_hd__a2bb2o_4
X_21596_ _15899_/A _21109_/B _21113_/C _21595_/X VGND VGND VPWR VPWR _21596_/X sky130_fd_sc_hd__a211o_4
X_24384_ _24361_/CLK _15942_/X HRESETn VGND VGND VPWR VPWR _22783_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20547_ _20545_/Y _20546_/Y _13515_/X VGND VGND VPWR VPWR _20547_/X sky130_fd_sc_hd__o21a_4
XFILLER_126_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23335_ _24750_/CLK _19437_/X VGND VGND VPWR VPWR _23335_/Q sky130_fd_sc_hd__dfxtp_4
X_20478_ _13508_/C _20474_/X _20477_/Y VGND VGND VPWR VPWR _20478_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24951__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23266_ _23242_/CLK _23266_/D VGND VGND VPWR VPWR _19633_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25005_ _25005_/CLK _13008_/X HRESETn VGND VGND VPWR VPWR _25005_/Q sky130_fd_sc_hd__dfrtp_4
X_22217_ _11529_/A _21106_/X VGND VGND VPWR VPWR _22510_/C sky130_fd_sc_hd__or2_4
XFILLER_105_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24269__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23197_ _23179_/CLK _19819_/X VGND VGND VPWR VPWR _19817_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__12125__A _24550_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16656__B1 _15501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12390__B1 _21104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22148_ _22148_/A VGND VGND VPWR VPWR _22148_/X sky130_fd_sc_hd__buf_2
XANTENNA__21438__A _21570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11964__A _11964_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14970_ _14964_/Y VGND VGND VPWR VPWR _15224_/A sky130_fd_sc_hd__buf_2
X_22079_ _21786_/A _22079_/B VGND VGND VPWR VPWR _22079_/X sky130_fd_sc_hd__or2_4
XFILLER_0_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13921_ _13921_/A VGND VGND VPWR VPWR _13934_/A sky130_fd_sc_hd__inv_2
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21401__B1 _13446_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16640_ _14713_/Y _16639_/X _16334_/X _16639_/X VGND VGND VPWR VPWR _24114_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17651__A _17651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13852_ _13852_/A _13849_/Y _13872_/C _13851_/X VGND VGND VPWR VPWR _13852_/X sky130_fd_sc_hd__or4_4
XFILLER_90_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_67_0_HCLK clkbuf_8_67_0_HCLK/A VGND VGND VPWR VPWR _24980_/CLK sky130_fd_sc_hd__clkbuf_1
X_12803_ _22779_/A VGND VGND VPWR VPWR _12803_/Y sky130_fd_sc_hd__inv_2
X_16571_ _14825_/Y _16570_/X _16141_/X _16570_/X VGND VGND VPWR VPWR _16571_/X sky130_fd_sc_hd__a2bb2o_4
X_13783_ _13761_/B VGND VGND VPWR VPWR _13783_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13642__B1 _13398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21704__A1 _21564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23833__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18310_ _18213_/D _18307_/B VGND VGND VPWR VPWR _18310_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22901__B1 _24054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15522_ _11630_/A VGND VGND VPWR VPWR _15522_/X sky130_fd_sc_hd__buf_2
XFILLER_128_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25057__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12734_ _12734_/A VGND VGND VPWR VPWR _12734_/Y sky130_fd_sc_hd__inv_2
X_19290_ _21827_/B _19284_/X _11844_/X _19289_/X VGND VGND VPWR VPWR _23388_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18241_ _18200_/Y _18240_/X VGND VGND VPWR VPWR _18257_/B sky130_fd_sc_hd__or2_4
X_15453_ _15453_/A VGND VGND VPWR VPWR _15453_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12665_ _12636_/X VGND VGND VPWR VPWR _13007_/B sky130_fd_sc_hd__inv_2
XFILLER_42_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16803__A1_N _24417_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _14384_/X _14399_/X _14402_/Y _14403_/X _13432_/A VGND VGND VPWR VPWR _24763_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _13665_/A VGND VGND VPWR VPWR _11616_/X sky130_fd_sc_hd__buf_2
X_18172_ _18172_/A _18172_/B _18172_/C _18172_/D VGND VGND VPWR VPWR _18172_/X sky130_fd_sc_hd__or4_4
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15384_ _15383_/Y _15381_/X _11607_/X _15381_/X VGND VGND VPWR VPWR _24592_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12596_ _12596_/A VGND VGND VPWR VPWR _12596_/Y sky130_fd_sc_hd__inv_2
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17123_ _17086_/A VGND VGND VPWR VPWR _17129_/A sky130_fd_sc_hd__buf_2
X_14335_ _23649_/Q VGND VGND VPWR VPWR _14335_/X sky130_fd_sc_hd__buf_2
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11547_ _11547_/A VGND VGND VPWR VPWR _11547_/Y sky130_fd_sc_hd__inv_2
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17054_ _17054_/A _17054_/B VGND VGND VPWR VPWR _17055_/B sky130_fd_sc_hd__or2_4
X_14266_ _13934_/A VGND VGND VPWR VPWR _14266_/X sky130_fd_sc_hd__buf_2
XANTENNA__24692__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16005_ _16005_/A VGND VGND VPWR VPWR _16005_/X sky130_fd_sc_hd__buf_2
X_13217_ _13146_/A _13217_/B VGND VGND VPWR VPWR _13218_/C sky130_fd_sc_hd__or2_4
XANTENNA__22432__A2 _20821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24621__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14197_ _14197_/A _14196_/X VGND VGND VPWR VPWR _14199_/B sky130_fd_sc_hd__or2_4
XANTENNA__19833__B1 _19832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13148_ _11743_/A _23340_/Q VGND VGND VPWR VPWR _13150_/B sky130_fd_sc_hd__or2_4
XFILLER_83_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13079_ _13166_/A _23597_/Q VGND VGND VPWR VPWR _13079_/X sky130_fd_sc_hd__or2_4
X_17956_ _17781_/A _17956_/B VGND VGND VPWR VPWR _17958_/B sky130_fd_sc_hd__or2_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16907_ _16824_/A _16907_/B VGND VGND VPWR VPWR _16907_/X sky130_fd_sc_hd__or2_4
X_17887_ _17887_/A _23417_/Q VGND VGND VPWR VPWR _17889_/B sky130_fd_sc_hd__or2_4
XFILLER_66_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19626_ _23269_/Q VGND VGND VPWR VPWR _21912_/B sky130_fd_sc_hd__inv_2
X_16838_ _16838_/A _16834_/X _16837_/X VGND VGND VPWR VPWR _16838_/X sky130_fd_sc_hd__or3_4
XFILLER_93_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16769_ _24083_/Q VGND VGND VPWR VPWR _16769_/Y sky130_fd_sc_hd__inv_2
X_19557_ _23293_/Q VGND VGND VPWR VPWR _21934_/B sky130_fd_sc_hd__inv_2
XANTENNA__13633__B1 _13632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18508_ _18508_/A VGND VGND VPWR VPWR _18509_/B sky130_fd_sc_hd__inv_2
X_19488_ _19487_/X VGND VGND VPWR VPWR _19488_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21811__A _20972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18439_ _18462_/A _18438_/X VGND VGND VPWR VPWR _18446_/A sky130_fd_sc_hd__or2_4
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21450_ _15281_/Y _11501_/X _24858_/Q _20758_/X VGND VGND VPWR VPWR _21450_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20401_ _20401_/A _20401_/B VGND VGND VPWR VPWR _20401_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_4_10_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_10_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_21381_ _14471_/X _21373_/X _21381_/C VGND VGND VPWR VPWR _21381_/X sky130_fd_sc_hd__or3_4
XANTENNA__22671__A2 _21896_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24709__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20332_ _20332_/A _20179_/B VGND VGND VPWR VPWR _20332_/Y sky130_fd_sc_hd__nand2_4
X_23120_ _23401_/CLK _20028_/X VGND VGND VPWR VPWR _20026_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__20682__B2 _20602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23051_ VGND VGND VPWR VPWR _23051_/HI sda_o_S5 sky130_fd_sc_hd__conb_1
X_20263_ _23764_/Q _20265_/B _20229_/X _20262_/X VGND VGND VPWR VPWR _20263_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24362__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22002_ _21245_/X _22002_/B _21999_/X _22002_/D VGND VGND VPWR VPWR _22002_/X sky130_fd_sc_hd__or4_4
XANTENNA__22361__B _21543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16638__B1 HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24023__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20194_ _20194_/A _20194_/B _20194_/C _20252_/A VGND VGND VPWR VPWR _20194_/X sky130_fd_sc_hd__or4_4
XFILLER_27_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18339__A1_N _16445_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23953_ _23949_/CLK _23953_/D HRESETn VGND VGND VPWR VPWR _22307_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_220_0_HCLK clkbuf_8_221_0_HCLK/A VGND VGND VPWR VPWR _23828_/CLK sky130_fd_sc_hd__clkbuf_1
X_22904_ _22900_/X _22904_/B _22902_/X _22903_/X VGND VGND VPWR VPWR _22904_/X sky130_fd_sc_hd__or4_4
XANTENNA__21705__B _21705_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23884_ _23885_/CLK _18116_/X HRESETn VGND VGND VPWR VPWR _18115_/A sky130_fd_sc_hd__dfrtp_4
X_22835_ _22835_/A VGND VGND VPWR VPWR _22835_/X sky130_fd_sc_hd__buf_2
XANTENNA__16087__A _16087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25150__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22766_ _16160_/A _22897_/B VGND VGND VPWR VPWR _22766_/X sky130_fd_sc_hd__or2_4
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24505_ _24502_/CLK _24505_/D HRESETn VGND VGND VPWR VPWR _24505_/Q sky130_fd_sc_hd__dfrtp_4
X_21717_ _21719_/A _21716_/X _16375_/Y _13618_/A VGND VGND VPWR VPWR _21717_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15377__B1 _11598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22697_ _22011_/X _22695_/X _21562_/X _22696_/X VGND VGND VPWR VPWR _22698_/A sky130_fd_sc_hd__o22a_4
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _25095_/Q _12449_/Y VGND VGND VPWR VPWR _12450_/X sky130_fd_sc_hd__or2_4
X_24436_ _24372_/CLK _24436_/D HRESETn VGND VGND VPWR VPWR _22126_/A sky130_fd_sc_hd__dfrtp_4
X_21648_ _21648_/A _20064_/X VGND VGND VPWR VPWR _21648_/X sky130_fd_sc_hd__and2_4
XFILLER_8_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12381_ _12379_/Y _21567_/A _25098_/Q _12380_/Y VGND VGND VPWR VPWR _12387_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22662__A2 _22536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24367_ _24361_/CLK _24367_/D HRESETn VGND VGND VPWR VPWR _24367_/Q sky130_fd_sc_hd__dfrtp_4
X_21579_ _21285_/B VGND VGND VPWR VPWR _22840_/A sky130_fd_sc_hd__buf_2
X_14120_ _14108_/A _14120_/B VGND VGND VPWR VPWR _14121_/C sky130_fd_sc_hd__or2_4
XFILLER_10_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23318_ _23332_/CLK _23318_/D VGND VGND VPWR VPWR _23318_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_125_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24298_ _24031_/CLK _24298_/D HRESETn VGND VGND VPWR VPWR _16195_/A sky130_fd_sc_hd__dfrtp_4
X_14051_ _14050_/Y _14048_/X _13665_/X _14048_/X VGND VGND VPWR VPWR _14051_/X sky130_fd_sc_hd__a2bb2o_4
X_23249_ _23249_/CLK _19681_/X VGND VGND VPWR VPWR _23249_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13002_ _12858_/X _13004_/B _13001_/Y VGND VGND VPWR VPWR _25008_/D sky130_fd_sc_hd__o21a_4
XANTENNA__21168__A _17651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24032__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22447__A2_N _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_30_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_61_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17810_ _17726_/A VGND VGND VPWR VPWR _17914_/A sky130_fd_sc_hd__buf_2
XFILLER_0_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18790_ _18798_/A VGND VGND VPWR VPWR _18790_/X sky130_fd_sc_hd__buf_2
XFILLER_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17741_ _17732_/A VGND VGND VPWR VPWR _17894_/A sky130_fd_sc_hd__buf_2
X_14953_ _24672_/Q VGND VGND VPWR VPWR _15136_/C sky130_fd_sc_hd__inv_2
XANTENNA__20800__A _20800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13904_ _13825_/X _13892_/X _13884_/X _13824_/X _13903_/X VGND VGND VPWR VPWR _13904_/X
+ sky130_fd_sc_hd__a32o_4
X_17672_ _17694_/A _18782_/A VGND VGND VPWR VPWR _17672_/X sky130_fd_sc_hd__or2_4
X_14884_ _14883_/Y _22312_/A _14883_/Y _22312_/A VGND VGND VPWR VPWR _14884_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16623_ _15619_/X _16597_/X _15743_/X _24124_/Q _16622_/X VGND VGND VPWR VPWR _16623_/X
+ sky130_fd_sc_hd__a32o_4
X_19411_ _19411_/A VGND VGND VPWR VPWR _19411_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16801__B1 _24415_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13835_ _13866_/B _13867_/A _13817_/X _13830_/X VGND VGND VPWR VPWR _13835_/X sky130_fd_sc_hd__or4_4
XFILLER_112_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16554_ _16553_/Y _16549_/X _16216_/X _16549_/X VGND VGND VPWR VPWR _16554_/X sky130_fd_sc_hd__a2bb2o_4
X_19342_ _19340_/Y _19341_/X _19227_/X _19341_/X VGND VGND VPWR VPWR _23369_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13766_ _13761_/B _13765_/Y _13782_/B _13766_/D VGND VGND VPWR VPWR _13767_/A sky130_fd_sc_hd__or4_4
X_15505_ HWDATA[12] VGND VGND VPWR VPWR _15505_/X sky130_fd_sc_hd__buf_2
XFILLER_31_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12717_ _12607_/Y _12714_/B VGND VGND VPWR VPWR _12717_/Y sky130_fd_sc_hd__nand2_4
X_19273_ _23393_/Q VGND VGND VPWR VPWR _19273_/Y sky130_fd_sc_hd__inv_2
X_16485_ _16485_/A VGND VGND VPWR VPWR _16485_/Y sky130_fd_sc_hd__inv_2
X_13697_ _23687_/Q VGND VGND VPWR VPWR _13697_/X sky130_fd_sc_hd__buf_2
X_18224_ _23876_/Q _18225_/B VGND VGND VPWR VPWR _18224_/X sky130_fd_sc_hd__or2_4
X_15436_ _14434_/A VGND VGND VPWR VPWR _15436_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12648_ _12648_/A VGND VGND VPWR VPWR _12648_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24873__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14040__B1 _13398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18155_ _18234_/A VGND VGND VPWR VPWR _18222_/B sky130_fd_sc_hd__inv_2
XFILLER_89_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15367_ _22487_/A _15366_/X _11581_/X _15366_/X VGND VGND VPWR VPWR _15367_/X sky130_fd_sc_hd__a2bb2o_4
X_12579_ _12579_/A VGND VGND VPWR VPWR _12579_/Y sky130_fd_sc_hd__inv_2
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17106_ _16982_/Y _17104_/X _17105_/Y VGND VGND VPWR VPWR _17106_/X sky130_fd_sc_hd__o21a_4
XFILLER_15_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14318_ _20177_/C _14317_/B _14329_/A _14317_/Y VGND VGND VPWR VPWR _14318_/X sky130_fd_sc_hd__a211o_4
X_18086_ _18086_/A VGND VGND VPWR VPWR _18086_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21861__B1 _14836_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15298_ _23761_/D _15297_/X VGND VGND VPWR VPWR _15298_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_112_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_225_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17037_ _24039_/Q VGND VGND VPWR VPWR _17043_/B sky130_fd_sc_hd__inv_2
X_14249_ _14248_/Y VGND VGND VPWR VPWR _14249_/X sky130_fd_sc_hd__buf_2
XFILLER_132_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22612__D _22611_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17293__B1 _11623_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16635__A3 HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18988_ _23494_/Q VGND VGND VPWR VPWR _22061_/B sky130_fd_sc_hd__inv_2
XANTENNA__19699__A1_N _19698_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17939_ _15729_/X _17923_/X _17938_/X _23928_/Q _15728_/A VGND VGND VPWR VPWR _17939_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__23755__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20950_ _20971_/A VGND VGND VPWR VPWR _22087_/A sky130_fd_sc_hd__buf_2
XANTENNA__17596__A1 _17490_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18793__B1 _18700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19609_ _23274_/Q VGND VGND VPWR VPWR _19609_/Y sky130_fd_sc_hd__inv_2
X_20881_ _20881_/A _20931_/A VGND VGND VPWR VPWR _20881_/Y sky130_fd_sc_hd__nand2_4
XPHY_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_50_0_HCLK clkbuf_8_51_0_HCLK/A VGND VGND VPWR VPWR _23990_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22620_ _24209_/Q _22580_/B VGND VGND VPWR VPWR _22620_/X sky130_fd_sc_hd__or2_4
XPHY_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22637__A _22637_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21541__A _13614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22551_ _22551_/A VGND VGND VPWR VPWR _22551_/X sky130_fd_sc_hd__buf_2
X_21502_ _21371_/A _21502_/B VGND VGND VPWR VPWR _21503_/C sky130_fd_sc_hd__or2_4
X_22482_ _22263_/X _22482_/B VGND VGND VPWR VPWR _22482_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__14031__B1 _13665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24221_ _24222_/CLK _16397_/X HRESETn VGND VGND VPWR VPWR _16389_/A sky130_fd_sc_hd__dfrtp_4
X_21433_ _24398_/Q _21292_/X _21107_/X _21432_/X VGND VGND VPWR VPWR _21433_/X sky130_fd_sc_hd__a211o_4
XFILLER_108_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24543__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21364_ _22806_/B _21362_/X _20745_/X _21363_/Y VGND VGND VPWR VPWR _21364_/X sky130_fd_sc_hd__a211o_4
XFILLER_107_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24152_ _24098_/CLK _16577_/X HRESETn VGND VGND VPWR VPWR _24152_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20315_ _18617_/B _20314_/Y _20315_/C VGND VGND VPWR VPWR _20315_/X sky130_fd_sc_hd__and3_4
X_23103_ _24962_/CLK _23103_/D VGND VGND VPWR VPWR _20069_/A sky130_fd_sc_hd__dfxtp_4
X_21295_ _24397_/Q _21292_/X _20744_/X _21294_/X VGND VGND VPWR VPWR _21296_/C sky130_fd_sc_hd__a211o_4
X_24083_ _24425_/CLK _16875_/X HRESETn VGND VGND VPWR VPWR _24083_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20246_ _20246_/A _20221_/B _14012_/Y _20232_/C VGND VGND VPWR VPWR _20246_/X sky130_fd_sc_hd__and4_4
X_23034_ _13622_/Y _23034_/B VGND VGND VPWR VPWR _23034_/Y sky130_fd_sc_hd__nor2_4
XFILLER_27_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_17_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20177_ _20177_/A _24780_/Q _20177_/C VGND VGND VPWR VPWR _20178_/A sky130_fd_sc_hd__or3_4
XFILLER_130_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16626__A3 HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12403__A _12508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24985_ _24776_/CLK _24985_/D HRESETn VGND VGND VPWR VPWR _11904_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21907__A1 _22223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11950_ _11949_/Y VGND VGND VPWR VPWR _11950_/X sky130_fd_sc_hd__buf_2
XFILLER_45_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23936_ _23486_/CLK _17664_/X HRESETn VGND VGND VPWR VPWR _13406_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_91_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15433__B _16475_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15598__B1 _11552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11881_ _11881_/A _11881_/B VGND VGND VPWR VPWR _11882_/B sky130_fd_sc_hd__and2_4
XFILLER_45_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23867_ _23859_/CLK _23867_/D HRESETn VGND VGND VPWR VPWR _23867_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13620_ _13611_/X _13619_/X VGND VGND VPWR VPWR _13620_/Y sky130_fd_sc_hd__nor2_4
XFILLER_44_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22818_ _21972_/X _22817_/X _22634_/X _24527_/Q _21187_/X VGND VGND VPWR VPWR _22818_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_77_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23798_ _23641_/CLK _20698_/X HRESETn VGND VGND VPWR VPWR _23798_/Q sky130_fd_sc_hd__dfrtp_4
X_13551_ _13550_/Y _13551_/B VGND VGND VPWR VPWR _13567_/B sky130_fd_sc_hd__or2_4
XFILLER_13_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22749_ _24213_/Q _22580_/B VGND VGND VPWR VPWR _22749_/X sky130_fd_sc_hd__or2_4
XANTENNA__16545__A HWDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12502_ _12502_/A _12409_/C VGND VGND VPWR VPWR _12502_/X sky130_fd_sc_hd__or2_4
XFILLER_12_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20894__A1 _22311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16270_ _16237_/A VGND VGND VPWR VPWR _16270_/X sky130_fd_sc_hd__buf_2
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13482_ _13480_/X VGND VGND VPWR VPWR _13482_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15221_ _15220_/X VGND VGND VPWR VPWR _24654_/D sky130_fd_sc_hd__inv_2
X_12433_ _12433_/A _12433_/B VGND VGND VPWR VPWR _12434_/C sky130_fd_sc_hd__or2_4
XFILLER_12_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24419_ _24425_/CLK _24419_/D HRESETn VGND VGND VPWR VPWR _15846_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24284__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15152_ _15152_/A VGND VGND VPWR VPWR _15156_/B sky130_fd_sc_hd__inv_2
X_12364_ _12465_/B _24481_/Q _12465_/B _24481_/Q VGND VGND VPWR VPWR _12364_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24213__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14103_ _13711_/X _20200_/A _14102_/X VGND VGND VPWR VPWR _14104_/A sky130_fd_sc_hd__o21a_4
X_15083_ _15059_/A _15059_/B _15016_/A _15080_/Y VGND VGND VPWR VPWR _15083_/X sky130_fd_sc_hd__a211o_4
X_19960_ _19960_/A VGND VGND VPWR VPWR _19960_/X sky130_fd_sc_hd__buf_2
X_12295_ _12293_/Y _12294_/X _12300_/C VGND VGND VPWR VPWR _12295_/X sky130_fd_sc_hd__and3_4
XFILLER_101_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14034_ _20209_/B VGND VGND VPWR VPWR _20221_/B sky130_fd_sc_hd__inv_2
X_18911_ _18910_/Y _18906_/X _18795_/X _18906_/X VGND VGND VPWR VPWR _18911_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19891_ _21784_/B _19885_/X _19821_/X _19890_/X VGND VGND VPWR VPWR _23172_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19803__A3 _13663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18842_ _23546_/Q VGND VGND VPWR VPWR _21506_/B sky130_fd_sc_hd__inv_2
XFILLER_79_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14089__B1 _13635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15985_ _15984_/Y _15979_/X _15890_/X _15979_/X VGND VGND VPWR VPWR _24367_/D sky130_fd_sc_hd__a2bb2o_4
X_18773_ _17860_/B VGND VGND VPWR VPWR _18773_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25072__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14936_ _14936_/A VGND VGND VPWR VPWR _14936_/Y sky130_fd_sc_hd__inv_2
X_17724_ _17815_/A _17724_/B _17724_/C VGND VGND VPWR VPWR _17739_/B sky130_fd_sc_hd__or3_4
XANTENNA__15624__A _15604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18000__A _11630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25001__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14867_ _14867_/A VGND VGND VPWR VPWR _15014_/A sky130_fd_sc_hd__buf_2
X_17655_ _15713_/X _16222_/C _15810_/X _17654_/X VGND VGND VPWR VPWR _17655_/X sky130_fd_sc_hd__a211o_4
XFILLER_24_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18935__A _18935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13144__A _13182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_37_0_HCLK clkbuf_6_18_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_75_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13818_ _13818_/A _13827_/A _13817_/X VGND VGND VPWR VPWR _13867_/C sky130_fd_sc_hd__or3_4
X_16606_ _16575_/A VGND VGND VPWR VPWR _16606_/X sky130_fd_sc_hd__buf_2
X_17586_ _17586_/A _17489_/X VGND VGND VPWR VPWR _17587_/B sky130_fd_sc_hd__or2_4
XFILLER_51_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14798_ _15035_/A _24143_/Q _15035_/A _24143_/Q VGND VGND VPWR VPWR _14798_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14261__B1 _14213_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16537_ _16537_/A VGND VGND VPWR VPWR _16537_/Y sky130_fd_sc_hd__inv_2
X_19325_ _13013_/B VGND VGND VPWR VPWR _19325_/Y sky130_fd_sc_hd__inv_2
X_13749_ _13769_/A _13769_/B _13764_/A VGND VGND VPWR VPWR _13757_/A sky130_fd_sc_hd__o21ai_4
XFILLER_91_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16455__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12395__A1_N _12408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16468_ _16467_/Y _16465_/X _16211_/X _16465_/X VGND VGND VPWR VPWR _16468_/X sky130_fd_sc_hd__a2bb2o_4
X_19256_ _25169_/Q VGND VGND VPWR VPWR _19256_/X sky130_fd_sc_hd__buf_2
X_15419_ _15411_/X _15415_/Y _15416_/X _20741_/B _15418_/X VGND VGND VPWR VPWR _15419_/X
+ sky130_fd_sc_hd__a32o_4
X_18207_ _18268_/A _18207_/B _18206_/X VGND VGND VPWR VPWR _18207_/X sky130_fd_sc_hd__or3_4
XANTENNA__11599__A _11599_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19187_ _19186_/Y _19182_/X _19120_/X _19175_/A VGND VGND VPWR VPWR _23423_/D sky130_fd_sc_hd__a2bb2o_4
X_16399_ _16398_/Y _16396_/X _16141_/X _16396_/X VGND VGND VPWR VPWR _24220_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_6_0_HCLK clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18138_ _16082_/Y _23861_/Q _16082_/Y _23861_/Q VGND VGND VPWR VPWR _18145_/A sky130_fd_sc_hd__a2bb2o_4
X_18069_ _11755_/Y _11729_/X _18075_/A VGND VGND VPWR VPWR _18069_/X sky130_fd_sc_hd__or3_4
X_20100_ _23092_/Q VGND VGND VPWR VPWR _21931_/B sky130_fd_sc_hd__inv_2
XANTENNA__12327__B1 _12412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21080_ _21079_/X VGND VGND VPWR VPWR _21080_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22920__A _22920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23936__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20031_ _23118_/Q VGND VGND VPWR VPWR _20947_/B sky130_fd_sc_hd__inv_2
XFILLER_99_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13038__B _13038_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15534__A _19442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24770_ _24769_/CLK _24770_/D HRESETn VGND VGND VPWR VPWR sda_oen_o_S4 sky130_fd_sc_hd__dfstp_4
X_21982_ _21178_/A _21980_/X _21981_/X _24508_/Q _16393_/D VGND VGND VPWR VPWR _21982_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17271__A2_N _17270_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23721_ _24180_/CLK _20533_/X HRESETn VGND VGND VPWR VPWR _13512_/C sky130_fd_sc_hd__dfrtp_4
X_20933_ _15426_/X _20932_/X _13546_/A _12062_/A VGND VGND VPWR VPWR _20933_/X sky130_fd_sc_hd__o22a_4
XPHY_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23652_ _23774_/CLK _23652_/D HRESETn VGND VGND VPWR VPWR _20158_/A sky130_fd_sc_hd__dfrtp_4
X_20864_ _20863_/X VGND VGND VPWR VPWR _20864_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24795__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15595__A3 _15477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22603_ _22129_/X _22602_/X _21994_/X _15862_/A _21995_/X VGND VGND VPWR VPWR _22603_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22865__A2 _22311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24724__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23583_ _23586_/CLK _18731_/X VGND VGND VPWR VPWR _17952_/B sky130_fd_sc_hd__dfxtp_4
X_20795_ _25190_/Q _20780_/X _20782_/X _20794_/X VGND VGND VPWR VPWR _20795_/X sky130_fd_sc_hd__a211o_4
XFILLER_23_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22534_ _22360_/X _22517_/X _22520_/X _22526_/X _22533_/X VGND VGND VPWR VPWR _22534_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_10_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14555__A1 _21257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22465_ _22299_/A _22464_/X VGND VGND VPWR VPWR _22465_/X sky130_fd_sc_hd__and2_4
XANTENNA__22814__B _20757_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24204_ _24201_/CLK _16440_/X HRESETn VGND VGND VPWR VPWR _16438_/A sky130_fd_sc_hd__dfrtp_4
X_21416_ _21040_/X _21413_/Y _22245_/A _21415_/X VGND VGND VPWR VPWR _21416_/X sky130_fd_sc_hd__a2bb2o_4
X_25184_ _25183_/CLK _11794_/X HRESETn VGND VGND VPWR VPWR _25184_/Q sky130_fd_sc_hd__dfrtp_4
X_22396_ _22396_/A _21978_/X VGND VGND VPWR VPWR _22398_/C sky130_fd_sc_hd__and2_4
XANTENNA__24808__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22533__C _22529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24135_ _24145_/CLK _16604_/X HRESETn VGND VGND VPWR VPWR _14831_/A sky130_fd_sc_hd__dfrtp_4
X_21347_ _21343_/X _21346_/X _21930_/A VGND VGND VPWR VPWR _21347_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15709__A _16216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12318__B1 _12416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12080_ _12079_/X _24570_/Q _12078_/Y _24570_/Q VGND VGND VPWR VPWR _12081_/D sky130_fd_sc_hd__a2bb2o_4
X_24066_ _24620_/CLK _24066_/D HRESETn VGND VGND VPWR VPWR _16771_/A sky130_fd_sc_hd__dfrtp_4
X_21278_ _16383_/A _21553_/A _20807_/X _21277_/X VGND VGND VPWR VPWR _21279_/C sky130_fd_sc_hd__a211o_4
XANTENNA__23677__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23017_ _24286_/Q _22859_/X _22338_/A VGND VGND VPWR VPWR _23017_/X sky130_fd_sc_hd__o21a_4
X_20229_ _20209_/A _15260_/A _20227_/X _20212_/D _20264_/B VGND VGND VPWR VPWR _20229_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15770_ HWDATA[20] VGND VGND VPWR VPWR _15770_/X sky130_fd_sc_hd__buf_2
X_12982_ _12982_/A VGND VGND VPWR VPWR _25015_/D sky130_fd_sc_hd__inv_2
X_24968_ _24968_/CLK _13490_/X HRESETn VGND VGND VPWR VPWR _13391_/B sky130_fd_sc_hd__dfstp_4
XFILLER_100_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14721_ _14876_/A VGND VGND VPWR VPWR _15035_/A sky130_fd_sc_hd__buf_2
XFILLER_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11933_ _11933_/A VGND VGND VPWR VPWR _11933_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23919_ _24937_/CLK _17991_/X HRESETn VGND VGND VPWR VPWR _22215_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_73_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20564__B1 _20562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24899_ _24902_/CLK _13915_/X HRESETn VGND VGND VPWR VPWR _24899_/Q sky130_fd_sc_hd__dfrtp_4
X_17440_ _17435_/X _17440_/B _17428_/C VGND VGND VPWR VPWR _17440_/X sky130_fd_sc_hd__and3_4
X_14652_ _23685_/D _14651_/Y _24628_/Q _23685_/D VGND VGND VPWR VPWR _14652_/X sky130_fd_sc_hd__a2bb2o_4
X_11864_ _21188_/A _11868_/A _11708_/B _13551_/B VGND VGND VPWR VPWR _11871_/C sky130_fd_sc_hd__o22a_4
XANTENNA__22277__A _22512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15586__A3 _15320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13603_ _13555_/X _13602_/Y _13553_/X _13586_/X _11687_/A VGND VGND VPWR VPWR _13603_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21181__A _21181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17371_ _17303_/Y _17348_/B VGND VGND VPWR VPWR _17371_/X sky130_fd_sc_hd__or2_4
X_14583_ _19946_/B VGND VGND VPWR VPWR _19123_/D sky130_fd_sc_hd__buf_2
XANTENNA__24465__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11795_ _11694_/X _11795_/B VGND VGND VPWR VPWR _11796_/B sky130_fd_sc_hd__or2_4
X_16322_ _16320_/Y _16321_/X _16153_/X _16321_/X VGND VGND VPWR VPWR _16322_/X sky130_fd_sc_hd__a2bb2o_4
X_19110_ _19108_/Y _19106_/X _19109_/X _19106_/X VGND VGND VPWR VPWR _23451_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13534_ _23737_/Q _13534_/B VGND VGND VPWR VPWR _20599_/A sky130_fd_sc_hd__or2_4
XFILLER_14_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19041_ _18743_/X VGND VGND VPWR VPWR _19041_/X sky130_fd_sc_hd__buf_2
X_16253_ _16228_/X _16234_/X _15600_/X _24278_/Q _16237_/X VGND VGND VPWR VPWR _16253_/X
+ sky130_fd_sc_hd__a32o_4
X_13465_ _21696_/A VGND VGND VPWR VPWR _13465_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15204_ _14883_/Y _15207_/B _15147_/X VGND VGND VPWR VPWR _15204_/Y sky130_fd_sc_hd__a21oi_4
X_12416_ _12416_/A _12415_/X VGND VGND VPWR VPWR _12417_/B sky130_fd_sc_hd__or2_4
X_16184_ _16196_/A VGND VGND VPWR VPWR _16184_/X sky130_fd_sc_hd__buf_2
X_13396_ _13396_/A VGND VGND VPWR VPWR SSn_S2 sky130_fd_sc_hd__inv_2
XFILLER_103_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15135_ _15135_/A VGND VGND VPWR VPWR _15135_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12347_ _12344_/A _12346_/A _12345_/X _12346_/Y VGND VGND VPWR VPWR _12351_/C sky130_fd_sc_hd__o22a_4
XANTENNA__15619__A _16624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12309__B1 _12417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15066_ _15078_/A _15061_/B VGND VGND VPWR VPWR _15079_/B sky130_fd_sc_hd__or2_4
X_19943_ _23151_/Q VGND VGND VPWR VPWR _19943_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12278_ _12261_/A _12278_/B _12277_/Y VGND VGND VPWR VPWR _12278_/X sky130_fd_sc_hd__and3_4
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14017_ _14016_/X VGND VGND VPWR VPWR _14197_/A sky130_fd_sc_hd__buf_2
XANTENNA__13139__A _13299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22241__B1 _25200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19874_ _21524_/B _19869_/X _19828_/X _19869_/X VGND VGND VPWR VPWR _23178_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22792__A1 _14850_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12147__A2_N _24571_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22792__B2 _22154_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18825_ _13258_/B VGND VGND VPWR VPWR _18825_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12978__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12777__A2_N _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18756_ _18756_/A VGND VGND VPWR VPWR _18756_/Y sky130_fd_sc_hd__inv_2
X_15968_ _24373_/Q VGND VGND VPWR VPWR _15968_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18748__B1 _18700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17707_ _17688_/X _17704_/X _17767_/A _23933_/Q _17705_/X VGND VGND VPWR VPWR _23933_/D
+ sky130_fd_sc_hd__a32o_4
X_14919_ _24679_/Q VGND VGND VPWR VPWR _15132_/A sky130_fd_sc_hd__inv_2
XFILLER_23_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15899_ _15899_/A VGND VGND VPWR VPWR _15899_/Y sky130_fd_sc_hd__inv_2
X_18687_ _13300_/B VGND VGND VPWR VPWR _18687_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17638_ _23940_/Q VGND VGND VPWR VPWR _17639_/A sky130_fd_sc_hd__buf_2
XFILLER_24_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17569_ _17568_/X VGND VGND VPWR VPWR _23958_/D sky130_fd_sc_hd__inv_2
XANTENNA__19173__B1 _19149_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19308_ _18739_/X VGND VGND VPWR VPWR _19308_/X sky130_fd_sc_hd__buf_2
X_20580_ _13532_/A _13532_/B _20579_/Y VGND VGND VPWR VPWR _20580_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24135__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_124_0_HCLK clkbuf_7_62_0_HCLK/X VGND VGND VPWR VPWR _23767_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_32_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_187_0_HCLK clkbuf_7_93_0_HCLK/X VGND VGND VPWR VPWR _25130_/CLK sky130_fd_sc_hd__clkbuf_1
X_19239_ _19238_/Y VGND VGND VPWR VPWR _19239_/X sky130_fd_sc_hd__buf_2
XFILLER_30_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22250_ _24477_/Q _22999_/B VGND VGND VPWR VPWR _22250_/X sky130_fd_sc_hd__or2_4
XFILLER_118_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21201_ _21500_/A _21201_/B _21200_/X VGND VGND VPWR VPWR _21201_/X sky130_fd_sc_hd__and3_4
XFILLER_69_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22181_ _21991_/X _22177_/X _20837_/X _22180_/Y VGND VGND VPWR VPWR _22181_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15529__A _15422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21132_ _21348_/A _21132_/B VGND VGND VPWR VPWR _21132_/X sky130_fd_sc_hd__or2_4
XANTENNA__23024__A2 _22285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22650__A _21050_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23770__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21063_ _21038_/X _21061_/X _21062_/X VGND VGND VPWR VPWR _21262_/A sky130_fd_sc_hd__o21a_4
XANTENNA__17744__A _17721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20014_ _20014_/A VGND VGND VPWR VPWR _20014_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11523__B2 _11521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18987__B1 _18964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24822_ _24823_/CLK _14205_/X HRESETn VGND VGND VPWR VPWR _24822_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24976__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14473__B1 _21396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24753_ _24757_/CLK _24753_/D HRESETn VGND VGND VPWR VPWR _13442_/A sky130_fd_sc_hd__dfrtp_4
X_21965_ _14488_/X _21964_/X _14494_/X VGND VGND VPWR VPWR _21965_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24905__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22809__B _20807_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ _23734_/CLK _20460_/Y HRESETn VGND VGND VPWR VPWR _13506_/C sky130_fd_sc_hd__dfrtp_4
X_20916_ _20911_/X _20915_/X _13441_/Y _20823_/X VGND VGND VPWR VPWR _20916_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24684_ _24264_/CLK _15091_/X HRESETn VGND VGND VPWR VPWR _24684_/Q sky130_fd_sc_hd__dfrtp_4
X_21896_ _22228_/A VGND VGND VPWR VPWR _21896_/X sky130_fd_sc_hd__buf_2
XPHY_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_20_0_HCLK clkbuf_7_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_20_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ _23641_/CLK _23635_/D HRESETn VGND VGND VPWR VPWR _20301_/A sky130_fd_sc_hd__dfrtp_4
X_20847_ _20847_/A VGND VGND VPWR VPWR _21093_/B sky130_fd_sc_hd__buf_2
XPHY_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21432__C _21432_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_83_0_HCLK clkbuf_7_83_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_83_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ HWDATA[15] VGND VGND VPWR VPWR _16087_/A sky130_fd_sc_hd__buf_2
XFILLER_126_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23566_ _24733_/CLK _23566_/D VGND VGND VPWR VPWR _18782_/A sky130_fd_sc_hd__dfxtp_4
X_20778_ _20778_/A _20777_/X VGND VGND VPWR VPWR _20778_/X sky130_fd_sc_hd__or2_4
XANTENNA__14851__A2_N _14850_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18911__B1 _18795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22517_ _22702_/A _22517_/B VGND VGND VPWR VPWR _22517_/X sky130_fd_sc_hd__and2_4
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23497_ _23128_/CLK _18983_/X VGND VGND VPWR VPWR _18981_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13250_ _13065_/X _13248_/X _13249_/X VGND VGND VPWR VPWR _13250_/X sky130_fd_sc_hd__and3_4
X_22448_ _21570_/X _22444_/X _22446_/X _20780_/X _22447_/X VGND VGND VPWR VPWR _22456_/C
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23858__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12201_ _12170_/A _12198_/X VGND VGND VPWR VPWR _12201_/X sky130_fd_sc_hd__or2_4
XFILLER_13_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15439__A _13454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13181_ _13271_/A VGND VGND VPWR VPWR _13222_/A sky130_fd_sc_hd__buf_2
X_25167_ _23898_/CLK _11872_/X HRESETn VGND VGND VPWR VPWR _25167_/Q sky130_fd_sc_hd__dfrtp_4
X_22379_ _21245_/X _22379_/B _22377_/X _22379_/D VGND VGND VPWR VPWR _22379_/X sky130_fd_sc_hd__or4_4
XFILLER_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12132_ _25115_/Q VGND VGND VPWR VPWR _12132_/Y sky130_fd_sc_hd__inv_2
X_24118_ _24112_/CLK _24118_/D HRESETn VGND VGND VPWR VPWR _24118_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16150__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22560__A _24306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25098_ _23716_/CLK _25098_/D HRESETn VGND VGND VPWR VPWR _25098_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21026__A1 _20908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12063_ _12062_/X VGND VGND VPWR VPWR _12063_/X sky130_fd_sc_hd__buf_2
X_16940_ _16940_/A VGND VGND VPWR VPWR _16951_/C sky130_fd_sc_hd__buf_2
X_24049_ _24049_/CLK _17093_/Y HRESETn VGND VGND VPWR VPWR _24049_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_46_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12711__B1 _12666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22774__A1 _22201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18978__B1 _18953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16871_ _16769_/Y _16874_/B VGND VGND VPWR VPWR _16875_/B sky130_fd_sc_hd__or2_4
X_18610_ _20288_/A _20283_/A VGND VGND VPWR VPWR _20289_/A sky130_fd_sc_hd__or2_4
X_15822_ _15414_/A _15821_/X VGND VGND VPWR VPWR _15822_/X sky130_fd_sc_hd__or2_4
X_19590_ _19590_/A VGND VGND VPWR VPWR _21223_/B sky130_fd_sc_hd__inv_2
XFILLER_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15753_ HWDATA[29] VGND VGND VPWR VPWR _15753_/X sky130_fd_sc_hd__buf_2
X_18541_ _18535_/A _18535_/B VGND VGND VPWR VPWR _18541_/Y sky130_fd_sc_hd__nand2_4
X_12965_ _12964_/X VGND VGND VPWR VPWR _12965_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14804__A2_N _24153_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24646__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11916_ _11903_/X _11916_/B _11916_/C _11916_/D VGND VGND VPWR VPWR _11916_/X sky130_fd_sc_hd__or4_4
X_14704_ _14703_/X _24118_/Q _14703_/X _24118_/Q VGND VGND VPWR VPWR _14704_/X sky130_fd_sc_hd__a2bb2o_4
X_15684_ _15657_/X VGND VGND VPWR VPWR _15684_/X sky130_fd_sc_hd__buf_2
X_18472_ _18472_/A _18472_/B VGND VGND VPWR VPWR _18474_/B sky130_fd_sc_hd__or2_4
XFILLER_73_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12896_ _12911_/A VGND VGND VPWR VPWR _12896_/X sky130_fd_sc_hd__buf_2
XFILLER_18_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14216__B1 _14094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14635_ _14634_/X VGND VGND VPWR VPWR _14655_/A sky130_fd_sc_hd__buf_2
X_17423_ _17423_/A _17423_/B _17422_/Y VGND VGND VPWR VPWR _17423_/X sky130_fd_sc_hd__and3_4
XFILLER_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11847_ _19610_/A VGND VGND VPWR VPWR _11847_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15964__B1 _11581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14767__B2 _24116_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14566_ _14564_/X _14565_/X _14561_/X VGND VGND VPWR VPWR _24737_/D sky130_fd_sc_hd__o21a_4
X_17354_ _17362_/A _17354_/B _17354_/C VGND VGND VPWR VPWR _17354_/X sky130_fd_sc_hd__and3_4
X_11778_ _11777_/X VGND VGND VPWR VPWR _11828_/B sky130_fd_sc_hd__inv_2
XFILLER_105_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17705__A1 _15712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18902__B1 _18901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13517_ _13516_/X VGND VGND VPWR VPWR _13517_/Y sky130_fd_sc_hd__inv_2
X_16305_ _16305_/A VGND VGND VPWR VPWR _16305_/X sky130_fd_sc_hd__buf_2
X_17285_ _11623_/Y _23982_/Q _25218_/Q _17340_/A VGND VGND VPWR VPWR _17290_/B sky130_fd_sc_hd__a2bb2o_4
X_14497_ _14453_/X _14462_/X _14497_/C _14497_/D VGND VGND VPWR VPWR _14497_/X sky130_fd_sc_hd__or4_4
XANTENNA__16733__A _22920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21550__A1_N _20235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16236_ _16240_/A VGND VGND VPWR VPWR _16237_/A sky130_fd_sc_hd__buf_2
X_19024_ _19024_/A VGND VGND VPWR VPWR _21374_/B sky130_fd_sc_hd__inv_2
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13448_ _13446_/A _13447_/A _13446_/Y _14374_/A VGND VGND VPWR VPWR _13448_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22309__A1_N _12508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16167_ _24309_/Q VGND VGND VPWR VPWR _16167_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13379_ _24978_/Q VGND VGND VPWR VPWR _13391_/A sky130_fd_sc_hd__inv_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15118_ _14966_/Y _15123_/A _15125_/A _15117_/X VGND VGND VPWR VPWR _15118_/X sky130_fd_sc_hd__or4_4
XFILLER_126_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23768__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16098_ _24335_/Q VGND VGND VPWR VPWR _16098_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15049_ _14878_/A _15123_/B VGND VGND VPWR VPWR _15049_/X sky130_fd_sc_hd__or2_4
X_19926_ _19925_/X VGND VGND VPWR VPWR _19926_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21568__A2 _21292_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21086__A _22014_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19857_ _21215_/B _19854_/X _19835_/X _19854_/X VGND VGND VPWR VPWR _23184_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18808_ _18807_/X VGND VGND VPWR VPWR _18809_/A sky130_fd_sc_hd__inv_2
XANTENNA__17641__B1 _17639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19788_ _23211_/Q VGND VGND VPWR VPWR _19788_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18739_ HWDATA[6] VGND VGND VPWR VPWR _18739_/X sky130_fd_sc_hd__buf_2
XANTENNA__24387__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21750_ _21751_/A _21251_/A VGND VGND VPWR VPWR _21750_/X sky130_fd_sc_hd__and2_4
XFILLER_58_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24316__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14207__B1 _13668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20701_ _20701_/A _14198_/X VGND VGND VPWR VPWR _20701_/X sky130_fd_sc_hd__and2_4
XFILLER_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15531__B _15531_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21681_ _21677_/A _19788_/Y VGND VGND VPWR VPWR _21681_/X sky130_fd_sc_hd__or2_4
XANTENNA__14758__B2 _24105_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14428__A _14428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23420_ _23596_/CLK _19197_/X VGND VGND VPWR VPWR _23420_/Q sky130_fd_sc_hd__dfxtp_4
X_20632_ _20635_/A _20627_/A _20631_/X VGND VGND VPWR VPWR _20632_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13430__A1 _13428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22645__A _24308_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19252__A2_N _19251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15707__B1 _24470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23351_ _23353_/CLK _23351_/D VGND VGND VPWR VPWR _19391_/A sky130_fd_sc_hd__dfxtp_4
X_20563_ _13525_/Y _13527_/B _13529_/B VGND VGND VPWR VPWR _20563_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16643__A _16643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22302_ _22302_/A VGND VGND VPWR VPWR _22302_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16380__B1 _15992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23282_ _23282_/CLK _19586_/X VGND VGND VPWR VPWR _19585_/A sky130_fd_sc_hd__dfxtp_4
X_20494_ _20499_/A VGND VGND VPWR VPWR _20495_/C sky130_fd_sc_hd__inv_2
XFILLER_30_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23951__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22083__C _22067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25021_ _25021_/CLK _25021_/D HRESETn VGND VGND VPWR VPWR _22527_/A sky130_fd_sc_hd__dfrtp_4
X_22233_ _22226_/X _22232_/X _16363_/Y _22228_/X VGND VGND VPWR VPWR _22233_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25175__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25104__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22164_ _22164_/A _22952_/B VGND VGND VPWR VPWR _22164_/X sky130_fd_sc_hd__or2_4
XFILLER_121_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21115_ _21112_/X _21867_/A VGND VGND VPWR VPWR _21127_/B sky130_fd_sc_hd__nor2_4
XFILLER_132_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16683__B2 _22307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22095_ _20946_/X _22095_/B VGND VGND VPWR VPWR _22095_/X sky130_fd_sc_hd__or2_4
XFILLER_82_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21046_ _22197_/A VGND VGND VPWR VPWR _21046_/X sky130_fd_sc_hd__buf_2
XFILLER_101_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24805_ _24823_/CLK _14254_/X HRESETn VGND VGND VPWR VPWR _24805_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_62_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22997_ _22997_/A _22997_/B _22990_/X _22996_/Y VGND VGND VPWR VPWR _22997_/X sky130_fd_sc_hd__or4_4
XFILLER_131_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12750_ _12647_/B _12741_/B VGND VGND VPWR VPWR _12751_/C sky130_fd_sc_hd__nand2_4
X_24736_ _23469_/CLK _14575_/X HRESETn VGND VGND VPWR VPWR _17674_/A sky130_fd_sc_hd__dfrtp_4
X_21948_ _21372_/A _21946_/X _21947_/X VGND VGND VPWR VPWR _21948_/X sky130_fd_sc_hd__and3_4
XANTENNA__16199__B1 _15982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21443__B _21097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24057__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11698_/C _11698_/D _11701_/C _11706_/A VGND VGND VPWR VPWR _11702_/B sky130_fd_sc_hd__and4_4
XFILLER_70_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12547_/A _12685_/B VGND VGND VPWR VPWR _12683_/B sky130_fd_sc_hd__or2_4
XANTENNA__15946__B1 _15765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24667_ _24671_/CLK _24667_/D HRESETn VGND VGND VPWR VPWR _24667_/Q sky130_fd_sc_hd__dfrtp_4
X_21879_ _21874_/X _21878_/X _13337_/A VGND VGND VPWR VPWR _21879_/X sky130_fd_sc_hd__o21a_4
XPHY_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14420_/A _14420_/B VGND VGND VPWR VPWR _14420_/X sky130_fd_sc_hd__or2_4
XPHY_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11628_/Y _11621_/X _11631_/X _11621_/X VGND VGND VPWR VPWR _25193_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23618_ _23618_/CLK _20157_/X HRESETn VGND VGND VPWR VPWR _23618_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24598_ _24596_/CLK _24598_/D HRESETn VGND VGND VPWR VPWR _24598_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22555__A _11961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14351_ _13811_/X _14350_/Y _13822_/X VGND VGND VPWR VPWR _14352_/C sky130_fd_sc_hd__o21a_4
XANTENNA__12794__A1_N _12793_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ HWDATA[20] VGND VGND VPWR VPWR _11563_/X sky130_fd_sc_hd__buf_2
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23549_ _23489_/CLK _18836_/X VGND VGND VPWR VPWR _23549_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13302_ _13238_/A _13302_/B _13302_/C VGND VGND VPWR VPWR _13303_/C sky130_fd_sc_hd__and3_4
XFILLER_7_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22274__B _22274_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17070_ _17070_/A _17070_/B VGND VGND VPWR VPWR _17070_/X sky130_fd_sc_hd__or2_4
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14282_ _24793_/Q VGND VGND VPWR VPWR _14282_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_170_0_HCLK clkbuf_7_85_0_HCLK/X VGND VGND VPWR VPWR _23308_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23692__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16021_ _16014_/B _16019_/X _16020_/Y VGND VGND VPWR VPWR _24357_/D sky130_fd_sc_hd__o21a_4
X_13233_ _13127_/A _20147_/A VGND VGND VPWR VPWR _13235_/B sky130_fd_sc_hd__or2_4
XANTENNA__15169__A _14950_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_27_0_HCLK clkbuf_8_27_0_HCLK/A VGND VGND VPWR VPWR _23411_/CLK sky130_fd_sc_hd__clkbuf_1
X_25219_ _23969_/CLK _11526_/X HRESETn VGND VGND VPWR VPWR _25219_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19864__A _19876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14921__B2 _14920_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23621__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22995__A1 _22429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13164_ _13073_/A _13158_/X _13164_/C VGND VGND VPWR VPWR _13164_/X sky130_fd_sc_hd__or3_4
XFILLER_100_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12115_ _12113_/A _24547_/Q _12265_/B _12114_/Y VGND VGND VPWR VPWR _12115_/X sky130_fd_sc_hd__o22a_4
XFILLER_124_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16674__B2 _16627_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13095_ _13090_/X _13092_/X _13094_/X VGND VGND VPWR VPWR _13095_/X sky130_fd_sc_hd__and3_4
X_17972_ _17705_/X _17971_/X _23926_/Q _17767_/A VGND VGND VPWR VPWR _23926_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24898__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22747__A1 _24148_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19711_ _11826_/A VGND VGND VPWR VPWR _19711_/X sky130_fd_sc_hd__buf_2
XANTENNA__16403__A1_N _16400_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12046_ _12045_/X VGND VGND VPWR VPWR _20697_/B sky130_fd_sc_hd__buf_2
X_16923_ _16923_/A _16942_/A VGND VGND VPWR VPWR _16924_/B sky130_fd_sc_hd__or2_4
XANTENNA__24827__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19642_ _20964_/B _19636_/X _19641_/X _19636_/A VGND VGND VPWR VPWR _19642_/X sky130_fd_sc_hd__a2bb2o_4
X_16854_ _16854_/A VGND VGND VPWR VPWR _16854_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15805_ _15439_/X VGND VGND VPWR VPWR _16222_/C sky130_fd_sc_hd__buf_2
X_19573_ _19573_/A VGND VGND VPWR VPWR _19573_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24480__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13997_ _13925_/A VGND VGND VPWR VPWR _13997_/Y sky130_fd_sc_hd__inv_2
X_16785_ _24412_/Q _16784_/Y _15896_/Y _24064_/Q VGND VGND VPWR VPWR _16785_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19376__B1 _19308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22449__B _20802_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18524_ _18427_/A _18523_/X VGND VGND VPWR VPWR _18545_/A sky130_fd_sc_hd__or2_4
XFILLER_92_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12948_ _12796_/Y _12947_/X VGND VGND VPWR VPWR _12949_/C sky130_fd_sc_hd__nand2_4
X_15736_ _15741_/B _16127_/A VGND VGND VPWR VPWR _15736_/X sky130_fd_sc_hd__or2_4
XFILLER_94_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18455_ _18412_/A _18453_/A VGND VGND VPWR VPWR _18455_/X sky130_fd_sc_hd__or2_4
XFILLER_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15937__B1 _11545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12879_ _22712_/A VGND VGND VPWR VPWR _12880_/C sky130_fd_sc_hd__inv_2
X_15667_ _12342_/Y _15666_/X _11525_/X _15666_/X VGND VGND VPWR VPWR _15667_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15674__A1_N _12332_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20930__B1 _20927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14758__A2_N _24105_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14248__A _15271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19128__B1 _19038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17406_ _17406_/A VGND VGND VPWR VPWR _17406_/Y sky130_fd_sc_hd__inv_2
X_14618_ _14618_/A _14618_/B _14617_/X VGND VGND VPWR VPWR _14619_/A sky130_fd_sc_hd__or3_4
XFILLER_18_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15598_ _12572_/Y _15593_/X _11552_/X _15593_/X VGND VGND VPWR VPWR _24526_/D sky130_fd_sc_hd__a2bb2o_4
X_18386_ _18380_/X _18383_/X _18384_/X _18385_/X VGND VGND VPWR VPWR _18386_/X sky130_fd_sc_hd__or4_4
X_14549_ _14543_/A VGND VGND VPWR VPWR _14549_/X sky130_fd_sc_hd__buf_2
X_17337_ _17330_/A _17329_/X _17331_/Y _17336_/X VGND VGND VPWR VPWR _17338_/A sky130_fd_sc_hd__a211o_4
XFILLER_53_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23709__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22184__B _22153_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17268_ _17261_/X _17263_/X _17265_/X _17267_/X VGND VGND VPWR VPWR _17269_/D sky130_fd_sc_hd__or4_4
XANTENNA__16362__B1 _16279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19007_ _23487_/Q VGND VGND VPWR VPWR _20990_/B sky130_fd_sc_hd__inv_2
X_16219_ _14218_/A VGND VGND VPWR VPWR _16219_/X sky130_fd_sc_hd__buf_2
X_17199_ _16369_/A VGND VGND VPWR VPWR _17199_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21809__A _20961_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19909_ _21962_/B _19906_/X _19818_/X _19906_/X VGND VGND VPWR VPWR _23165_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24568__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13327__A _16301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22920_ _22920_/A _23004_/A VGND VGND VPWR VPWR _22920_/X sky130_fd_sc_hd__and2_4
XFILLER_29_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21544__A _21544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13046__B _23598_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22851_ _22919_/A _22851_/B _22842_/X _22851_/D VGND VGND VPWR VPWR _22851_/X sky130_fd_sc_hd__or4_4
XANTENNA__19367__B1 _19366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21802_ _23976_/Q _20066_/Y _21799_/X _21801_/X VGND VGND VPWR VPWR _21802_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21263__B _21408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24150__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22782_ _22782_/A _22429_/B VGND VGND VPWR VPWR _22782_/X sky130_fd_sc_hd__or2_4
XFILLER_36_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21713__A2 _21707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24521_ _24521_/CLK _15608_/X HRESETn VGND VGND VPWR VPWR _24521_/Q sky130_fd_sc_hd__dfrtp_4
X_21733_ _21733_/A _21716_/B VGND VGND VPWR VPWR _21737_/A sky130_fd_sc_hd__and2_4
XFILLER_101_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18853__A _18852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24452_ _24459_/CLK _15764_/X HRESETn VGND VGND VPWR VPWR _24452_/Q sky130_fd_sc_hd__dfrtp_4
X_21664_ _21677_/A _18840_/Y VGND VGND VPWR VPWR _21664_/X sky130_fd_sc_hd__or2_4
XFILLER_40_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23403_ _23939_/CLK _19247_/X VGND VGND VPWR VPWR _19246_/A sky130_fd_sc_hd__dfxtp_4
X_20615_ _13535_/C _20611_/X _20614_/Y VGND VGND VPWR VPWR _20615_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_138_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24383_ _24385_/CLK _24383_/D HRESETn VGND VGND VPWR VPWR _22763_/A sky130_fd_sc_hd__dfrtp_4
X_21595_ _24293_/Q _20931_/A VGND VGND VPWR VPWR _21595_/X sky130_fd_sc_hd__and2_4
XFILLER_137_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16373__A _16373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23334_ _23308_/CLK _23334_/D VGND VGND VPWR VPWR _23334_/Q sky130_fd_sc_hd__dfxtp_4
X_20546_ _20542_/X VGND VGND VPWR VPWR _20546_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16353__B1 _15369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_243_0_HCLK clkbuf_8_243_0_HCLK/A VGND VGND VPWR VPWR _24104_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22426__B1 _20801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23265_ _23249_/CLK _23265_/D VGND VGND VPWR VPWR _23265_/Q sky130_fd_sc_hd__dfxtp_4
X_20477_ _13509_/C VGND VGND VPWR VPWR _20477_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25004_ _24944_/CLK _25004_/D HRESETn VGND VGND VPWR VPWR _13009_/A sky130_fd_sc_hd__dfrtp_4
X_22216_ _20918_/X _22214_/X _20903_/X _22215_/Y VGND VGND VPWR VPWR _22216_/X sky130_fd_sc_hd__o22a_4
X_23196_ _23154_/CLK _23196_/D VGND VGND VPWR VPWR _19820_/A sky130_fd_sc_hd__dfxtp_4
X_22147_ _22147_/A VGND VGND VPWR VPWR _22147_/X sky130_fd_sc_hd__buf_2
XFILLER_133_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24991__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22078_ _21760_/X _19508_/Y VGND VGND VPWR VPWR _22078_/X sky130_fd_sc_hd__or2_4
XFILLER_86_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24920__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13920_ _23694_/Q _13905_/A _13900_/X _13815_/X _13886_/X VGND VGND VPWR VPWR _13920_/X
+ sky130_fd_sc_hd__a32o_4
X_21029_ _20814_/X VGND VGND VPWR VPWR _21029_/X sky130_fd_sc_hd__buf_2
XFILLER_120_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21401__B2 _21400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24238__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_5_12_0_HCLK_A clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13851_ _13829_/X _13851_/B VGND VGND VPWR VPWR _13851_/X sky130_fd_sc_hd__or2_4
XANTENNA__19358__B1 _19221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12802_ _22778_/A VGND VGND VPWR VPWR _12802_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15452__A _14436_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13782_ _13764_/A _13782_/B _13780_/B VGND VGND VPWR VPWR _13787_/A sky130_fd_sc_hd__or3_4
X_16570_ _16570_/A VGND VGND VPWR VPWR _16570_/X sky130_fd_sc_hd__buf_2
XFILLER_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21704__A2 _21693_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12733_ _12728_/A _12728_/B _12730_/B _12666_/X VGND VGND VPWR VPWR _12734_/A sky130_fd_sc_hd__a211o_4
X_15521_ _15503_/X _15504_/X _15520_/X _24549_/Q _15466_/A VGND VGND VPWR VPWR _24549_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19859__A _19859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24719_ _24723_/CLK _14675_/X HRESETn VGND VGND VPWR VPWR _24719_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18763__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15452_ _14436_/B _15452_/B VGND VGND VPWR VPWR _15452_/Y sky130_fd_sc_hd__nor2_4
X_18240_ _18263_/A _18263_/B _18240_/C _18207_/X VGND VGND VPWR VPWR _18240_/X sky130_fd_sc_hd__or4_4
X_12664_ _12641_/X _12663_/X VGND VGND VPWR VPWR _12664_/X sky130_fd_sc_hd__or2_4
XFILLER_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21901__B _21720_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16592__B1 _16266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22285__A _21020_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23873__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14403_/A VGND VGND VPWR VPWR _14403_/X sky130_fd_sc_hd__buf_2
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ HWDATA[6] VGND VGND VPWR VPWR _13665_/A sky130_fd_sc_hd__buf_2
XANTENNA__22716__C _22716_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25097__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_53_0_HCLK clkbuf_6_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_53_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15383_ _24592_/Q VGND VGND VPWR VPWR _15383_/Y sky130_fd_sc_hd__inv_2
X_18171_ _16089_/Y _23859_/Q _16089_/Y _23859_/Q VGND VGND VPWR VPWR _18172_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ _24503_/Q VGND VGND VPWR VPWR _12595_/Y sky130_fd_sc_hd__inv_2
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23802__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14334_ _14329_/A _14333_/X _24790_/Q _14331_/X VGND VGND VPWR VPWR _14334_/X sky130_fd_sc_hd__o22a_4
X_17122_ _17122_/A VGND VGND VPWR VPWR _17122_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25026__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11546_ _11544_/Y _11542_/X _11545_/X _11542_/X VGND VGND VPWR VPWR _11546_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16344__B1 _16266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19712__A2_N _19710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17053_ _17053_/A _17086_/A VGND VGND VPWR VPWR _17054_/B sky130_fd_sc_hd__and2_4
X_14265_ _14264_/Y _14260_/X _14218_/X _14248_/Y VGND VGND VPWR VPWR _14265_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22417__B1 _22404_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12316__A _24477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16004_ _16003_/Y _14435_/B VGND VGND VPWR VPWR _16005_/A sky130_fd_sc_hd__or2_4
XANTENNA__22732__B _22953_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13216_ _13092_/A _13216_/B VGND VGND VPWR VPWR _13218_/B sky130_fd_sc_hd__or2_4
X_14196_ _16231_/A _21072_/A VGND VGND VPWR VPWR _14196_/X sky130_fd_sc_hd__or2_4
X_13147_ _13102_/X _13144_/X _13147_/C VGND VGND VPWR VPWR _13147_/X sky130_fd_sc_hd__and3_4
XANTENNA__21640__B2 _22616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13078_ _13078_/A VGND VGND VPWR VPWR _13166_/A sky130_fd_sc_hd__buf_2
X_17955_ _17955_/A _17947_/X _17955_/C VGND VGND VPWR VPWR _17955_/X sky130_fd_sc_hd__and3_4
XFILLER_65_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24661__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12133__B2 _24558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12029_ _12016_/B VGND VGND VPWR VPWR _12029_/Y sky130_fd_sc_hd__inv_2
X_16906_ _16893_/X VGND VGND VPWR VPWR _16907_/B sky130_fd_sc_hd__inv_2
XFILLER_66_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13147__A _13102_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17886_ _17780_/A _17886_/B _17886_/C VGND VGND VPWR VPWR _17890_/B sky130_fd_sc_hd__and3_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19625_ _22087_/B _19624_/X _19597_/X _19624_/X VGND VGND VPWR VPWR _23270_/D sky130_fd_sc_hd__a2bb2o_4
X_16837_ _16923_/A _16922_/A _16921_/C _16837_/D VGND VGND VPWR VPWR _16837_/X sky130_fd_sc_hd__or4_4
XANTENNA__11892__B1 _11890_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19556_ _22109_/B _19555_/X _11835_/X _19555_/X VGND VGND VPWR VPWR _23294_/D sky130_fd_sc_hd__a2bb2o_4
X_16768_ _24403_/Q _24067_/Q _15887_/Y _16935_/A VGND VGND VPWR VPWR _16773_/B sky130_fd_sc_hd__o22a_4
XFILLER_34_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18507_ _18486_/B _18507_/B VGND VGND VPWR VPWR _18508_/A sky130_fd_sc_hd__or2_4
X_15719_ _15713_/X VGND VGND VPWR VPWR _15720_/A sky130_fd_sc_hd__inv_2
XANTENNA__11644__B1 _11643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19487_ _14540_/X _19883_/B _19883_/C VGND VGND VPWR VPWR _19487_/X sky130_fd_sc_hd__or3_4
X_16699_ _16699_/A VGND VGND VPWR VPWR _16700_/A sky130_fd_sc_hd__inv_2
X_18438_ _18438_/A _18438_/B VGND VGND VPWR VPWR _18438_/X sky130_fd_sc_hd__or2_4
XFILLER_22_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22195__A _20753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18369_ _24209_/Q _23832_/Q _16425_/Y _18434_/C VGND VGND VPWR VPWR _18369_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16193__A _16193_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14706__A _24698_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20400_ _15270_/Y _17187_/X _17170_/Y _17184_/Y VGND VGND VPWR VPWR _20401_/B sky130_fd_sc_hd__o22a_4
XANTENNA__13610__A _16301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21380_ _21376_/X _21379_/X _21242_/X VGND VGND VPWR VPWR _21381_/C sky130_fd_sc_hd__o21a_4
XANTENNA__16335__B1 _16334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22923__A _22982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20331_ _20331_/A _20179_/B VGND VGND VPWR VPWR _20333_/B sky130_fd_sc_hd__or2_4
XFILLER_135_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_10_0_HCLK clkbuf_7_5_0_HCLK/X VGND VGND VPWR VPWR _23293_/CLK sky130_fd_sc_hd__clkbuf_1
X_23050_ VGND VGND VPWR VPWR _23050_/HI sda_o_S4 sky130_fd_sc_hd__conb_1
X_20262_ _15250_/A _20212_/B _23771_/Q _20264_/A VGND VGND VPWR VPWR _20262_/X sky130_fd_sc_hd__and4_4
XANTENNA__24749__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22001_ _12408_/C _22259_/A _25011_/Q _21051_/X VGND VGND VPWR VPWR _22002_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_73_0_HCLK clkbuf_7_36_0_HCLK/X VGND VGND VPWR VPWR _25141_/CLK sky130_fd_sc_hd__clkbuf_1
X_20193_ _20193_/A _20189_/B _20193_/C _20192_/X VGND VGND VPWR VPWR _20252_/A sky130_fd_sc_hd__and4_4
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13321__B1 _24996_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23952_ _23972_/CLK _17597_/Y HRESETn VGND VGND VPWR VPWR _22256_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_29_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24331__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21395__B1 _21242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22903_ _20534_/Y _20926_/X _13540_/A _22657_/X VGND VGND VPWR VPWR _22903_/X sky130_fd_sc_hd__a2bb2o_4
X_23883_ _23885_/CLK _18119_/X HRESETn VGND VGND VPWR VPWR _23883_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_44_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22834_ _24315_/Q _22834_/B VGND VGND VPWR VPWR _22834_/X sky130_fd_sc_hd__or2_4
XFILLER_129_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18012__B1 _16671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22765_ _22764_/X VGND VGND VPWR VPWR _22765_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24504_ _25009_/CLK _24504_/D HRESETn VGND VGND VPWR VPWR _12585_/A sky130_fd_sc_hd__dfrtp_4
X_21716_ _21716_/A _21716_/B VGND VGND VPWR VPWR _21716_/X sky130_fd_sc_hd__and2_4
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16574__B1 _24153_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22696_ _22696_/A _22587_/B VGND VGND VPWR VPWR _22696_/X sky130_fd_sc_hd__and2_4
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17199__A _16369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25190__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24435_ _24435_/CLK _15794_/X HRESETn VGND VGND VPWR VPWR _21980_/A sky130_fd_sc_hd__dfrtp_4
X_21647_ _21648_/A _20064_/X _18089_/Y _23104_/Q VGND VGND VPWR VPWR _21647_/X sky130_fd_sc_hd__o22a_4
XFILLER_123_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12380_ _24495_/Q VGND VGND VPWR VPWR _12380_/Y sky130_fd_sc_hd__inv_2
X_24366_ _24590_/CLK _24366_/D HRESETn VGND VGND VPWR VPWR _24366_/Q sky130_fd_sc_hd__dfrtp_4
X_21578_ _21570_/X _21572_/X _21574_/X _20800_/X _21577_/X VGND VGND VPWR VPWR _21602_/C
+ sky130_fd_sc_hd__a32o_4
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22833__A _22249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23317_ _23313_/CLK _19492_/X VGND VGND VPWR VPWR _19491_/A sky130_fd_sc_hd__dfxtp_4
X_20529_ _20527_/Y _20524_/Y _20528_/X VGND VGND VPWR VPWR _20529_/X sky130_fd_sc_hd__o21a_4
XFILLER_123_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24297_ _24319_/CLK _24297_/D HRESETn VGND VGND VPWR VPWR _16198_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_10_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14050_ _14050_/A VGND VGND VPWR VPWR _14050_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23248_ _23249_/CLK _19683_/X VGND VGND VPWR VPWR _19682_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_49_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13001_ _12858_/X _13004_/B _12896_/X VGND VGND VPWR VPWR _13001_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24419__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23179_ _23179_/CLK _23179_/D VGND VGND VPWR VPWR _19871_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_67_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17740_ _14563_/A VGND VGND VPWR VPWR _17898_/A sky130_fd_sc_hd__buf_2
X_14952_ _14945_/X _14947_/X _14949_/X _14951_/X VGND VGND VPWR VPWR _14973_/B sky130_fd_sc_hd__or4_4
XFILLER_130_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24072__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13903_ _13886_/X VGND VGND VPWR VPWR _13903_/X sky130_fd_sc_hd__buf_2
XANTENNA__18251__B1 _18228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17671_ _17697_/A _17671_/B VGND VGND VPWR VPWR _17673_/B sky130_fd_sc_hd__or2_4
XANTENNA__24001__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14883_ _24661_/Q VGND VGND VPWR VPWR _14883_/Y sky130_fd_sc_hd__inv_2
X_19410_ _19408_/Y _19409_/X _19387_/X _19409_/X VGND VGND VPWR VPWR _23345_/D sky130_fd_sc_hd__a2bb2o_4
X_16622_ _16627_/A VGND VGND VPWR VPWR _16622_/X sky130_fd_sc_hd__buf_2
XFILLER_21_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13834_ _13828_/A VGND VGND VPWR VPWR _13866_/B sky130_fd_sc_hd__buf_2
XFILLER_1_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19341_ _19327_/Y VGND VGND VPWR VPWR _19341_/X sky130_fd_sc_hd__buf_2
XFILLER_56_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18003__B1 _16617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13765_ _13764_/X _13761_/A VGND VGND VPWR VPWR _13765_/Y sky130_fd_sc_hd__nand2_4
X_16553_ _16553_/A VGND VGND VPWR VPWR _16553_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15504_ _15460_/X VGND VGND VPWR VPWR _15504_/X sky130_fd_sc_hd__buf_2
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15910__A _15916_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12716_ _12716_/A _12716_/B _12715_/Y VGND VGND VPWR VPWR _25055_/D sky130_fd_sc_hd__and3_4
X_19272_ _19271_/Y _19266_/X _19201_/X _19266_/X VGND VGND VPWR VPWR _19272_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25207__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13696_ _13678_/X _13695_/X _14081_/A _13693_/X VGND VGND VPWR VPWR _13696_/X sky130_fd_sc_hd__o22a_4
X_16484_ _16483_/Y _16481_/X _16243_/X _16481_/X VGND VGND VPWR VPWR _24187_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16724__A2_N _22376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18223_ _18223_/A _18223_/B VGND VGND VPWR VPWR _18225_/B sky130_fd_sc_hd__nor2_4
X_12647_ _12581_/Y _12647_/B _12647_/C _12739_/A VGND VGND VPWR VPWR _12652_/A sky130_fd_sc_hd__or4_4
X_15435_ _15435_/A VGND VGND VPWR VPWR _15438_/A sky130_fd_sc_hd__buf_2
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14526__A _14521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15366_ _15358_/X VGND VGND VPWR VPWR _15366_/X sky130_fd_sc_hd__buf_2
X_18154_ _18154_/A _18149_/X _18151_/X _18153_/X VGND VGND VPWR VPWR _18154_/X sky130_fd_sc_hd__or4_4
XANTENNA__16317__B1 _11536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12578_ _25066_/Q VGND VGND VPWR VPWR _12578_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17105_ _16982_/Y _17104_/X _17057_/X VGND VGND VPWR VPWR _17105_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11529_ _11529_/A VGND VGND VPWR VPWR _22992_/B sky130_fd_sc_hd__buf_2
X_14317_ _20177_/C _14317_/B VGND VGND VPWR VPWR _14317_/Y sky130_fd_sc_hd__nor2_4
XFILLER_129_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17837__A _17742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15297_ _15295_/A _15294_/Y _15296_/Y _14367_/Y VGND VGND VPWR VPWR _15297_/X sky130_fd_sc_hd__a211o_4
X_18085_ _18085_/A _18080_/A VGND VGND VPWR VPWR _18085_/X sky130_fd_sc_hd__and2_4
XANTENNA__21861__B2 _20757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14248_ _15271_/A _18633_/A VGND VGND VPWR VPWR _14248_/Y sky130_fd_sc_hd__nor2_4
X_17036_ _24040_/Q VGND VGND VPWR VPWR _17128_/A sky130_fd_sc_hd__inv_2
XANTENNA__24842__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14179_ _24830_/Q _14171_/X _24829_/Q _14176_/X VGND VGND VPWR VPWR _14179_/X sky130_fd_sc_hd__o22a_4
XFILLER_113_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18987_ _18986_/Y _18982_/X _18964_/X _18982_/A VGND VGND VPWR VPWR _18987_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17572__A _22473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17938_ _16022_/Y _17938_/B _17937_/X VGND VGND VPWR VPWR _17938_/X sky130_fd_sc_hd__and3_4
XFILLER_22_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11865__B1 _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17869_ _17961_/A _17869_/B _17869_/C VGND VGND VPWR VPWR _17873_/B sky130_fd_sc_hd__and3_4
X_19608_ _19606_/Y _19604_/X _19607_/X _19604_/X VGND VGND VPWR VPWR _19608_/X sky130_fd_sc_hd__a2bb2o_4
X_20880_ _20880_/A _11725_/X VGND VGND VPWR VPWR _20880_/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23795__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19539_ _19533_/Y VGND VGND VPWR VPWR _19539_/X sky130_fd_sc_hd__buf_2
XANTENNA__11617__B1 _11616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22877__B1 _22351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23724__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15820__A _22933_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22550_ _14838_/Y _22537_/X _14933_/Y _22549_/X VGND VGND VPWR VPWR _22550_/X sky130_fd_sc_hd__o22a_4
X_21501_ _21392_/A _21501_/B VGND VGND VPWR VPWR _21503_/B sky130_fd_sc_hd__or2_4
XFILLER_37_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22481_ _22225_/X _22478_/X _22231_/X _22480_/X VGND VGND VPWR VPWR _22482_/B sky130_fd_sc_hd__o22a_4
XFILLER_22_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24220_ _24225_/CLK _24220_/D HRESETn VGND VGND VPWR VPWR _16398_/A sky130_fd_sc_hd__dfrtp_4
X_21432_ _21432_/A _21431_/X _21432_/C VGND VGND VPWR VPWR _21432_/X sky130_fd_sc_hd__and3_4
XFILLER_108_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24151_ _24264_/CLK _24151_/D HRESETn VGND VGND VPWR VPWR _14859_/A sky130_fd_sc_hd__dfrtp_4
X_21363_ _21363_/A _11986_/X VGND VGND VPWR VPWR _21363_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__17747__A _17742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23102_ _23925_/CLK _20073_/X VGND VGND VPWR VPWR _20072_/A sky130_fd_sc_hd__dfxtp_4
X_20314_ _18616_/A _18616_/B VGND VGND VPWR VPWR _20314_/Y sky130_fd_sc_hd__nand2_4
X_24082_ _24079_/CLK _24082_/D HRESETn VGND VGND VPWR VPWR _16821_/A sky130_fd_sc_hd__dfrtp_4
X_21294_ _21432_/A _21293_/X _21432_/C VGND VGND VPWR VPWR _21294_/X sky130_fd_sc_hd__and3_4
XANTENNA__24583__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11795__A _11694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23033_ _13637_/Y _14428_/A _24942_/Q _20919_/A VGND VGND VPWR VPWR _23033_/X sky130_fd_sc_hd__a2bb2o_4
X_20245_ _20245_/A _20204_/X _20200_/A VGND VGND VPWR VPWR _20245_/X sky130_fd_sc_hd__and3_4
XFILLER_103_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24512__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20176_ _20234_/B VGND VGND VPWR VPWR _20179_/B sky130_fd_sc_hd__buf_2
XFILLER_76_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20901__A _22587_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12403__B _12403_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17482__A _17482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21716__B _21716_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24984_ _24984_/CLK _13367_/X HRESETn VGND VGND VPWR VPWR _11880_/A sky130_fd_sc_hd__dfrtp_4
X_23935_ _23486_/CLK _17668_/X HRESETn VGND VGND VPWR VPWR _13406_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15047__B1 _15027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11880_ _11880_/A VGND VGND VPWR VPWR _22006_/A sky130_fd_sc_hd__inv_2
X_23866_ _23762_/CLK _23866_/D HRESETn VGND VGND VPWR VPWR _23866_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11608__B1 _11607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22817_ _24454_/Q _22703_/B VGND VGND VPWR VPWR _22817_/X sky130_fd_sc_hd__or2_4
X_23797_ _23789_/CLK _20697_/X HRESETn VGND VGND VPWR VPWR _12016_/A sky130_fd_sc_hd__dfrtp_4
X_13550_ _23904_/Q VGND VGND VPWR VPWR _13550_/Y sky130_fd_sc_hd__inv_2
X_22748_ _22691_/A _22745_/X _22748_/C VGND VGND VPWR VPWR _22775_/A sky130_fd_sc_hd__and3_4
XANTENNA__16547__B1 _16546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12501_ _12500_/X VGND VGND VPWR VPWR _25082_/D sky130_fd_sc_hd__inv_2
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13481_ _13464_/X _13470_/B VGND VGND VPWR VPWR _13481_/X sky130_fd_sc_hd__or2_4
X_22679_ _12382_/A _22957_/B VGND VGND VPWR VPWR _22679_/X sky130_fd_sc_hd__and2_4
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15220_ _15197_/A _15197_/B _15218_/B _15147_/X VGND VGND VPWR VPWR _15220_/X sky130_fd_sc_hd__a211o_4
XANTENNA__13250__A _13065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12432_ _12432_/A _12432_/B VGND VGND VPWR VPWR _12434_/B sky130_fd_sc_hd__or2_4
X_24418_ _24425_/CLK _15850_/X HRESETn VGND VGND VPWR VPWR _15849_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22563__A _20814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15151_ _15154_/A _15146_/X _15151_/C VGND VGND VPWR VPWR _24674_/D sky130_fd_sc_hd__and3_4
X_12363_ _12411_/B VGND VGND VPWR VPWR _12465_/B sky130_fd_sc_hd__buf_2
X_24349_ _24349_/CLK _16062_/X HRESETn VGND VGND VPWR VPWR _16061_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14102_ _14072_/A _23658_/Q VGND VGND VPWR VPWR _14102_/X sky130_fd_sc_hd__or2_4
XANTENNA__22282__B _22281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15082_ _15057_/X _15061_/B _15081_/X VGND VGND VPWR VPWR _15082_/X sky130_fd_sc_hd__and3_4
XANTENNA__21179__A _21179_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12294_ _12265_/A _12293_/B VGND VGND VPWR VPWR _12294_/X sky130_fd_sc_hd__or2_4
XFILLER_4_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12336__A1 _25077_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14033_ _20246_/A _14026_/X _13668_/X _14028_/X VGND VGND VPWR VPWR _14033_/X sky130_fd_sc_hd__a2bb2o_4
X_18910_ _17868_/B VGND VGND VPWR VPWR _18910_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19890_ _19897_/A VGND VGND VPWR VPWR _19890_/X sky130_fd_sc_hd__buf_2
XANTENNA__24253__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18841_ _18840_/Y _18838_/X _15554_/X _18838_/X VGND VGND VPWR VPWR _18841_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18772_ _18771_/Y _18769_/X _18700_/X _18769_/X VGND VGND VPWR VPWR _23571_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15984_ _24367_/Q VGND VGND VPWR VPWR _15984_/Y sky130_fd_sc_hd__inv_2
X_17723_ _17716_/X _17719_/X _17723_/C VGND VGND VPWR VPWR _17724_/C sky130_fd_sc_hd__and3_4
XANTENNA__22020__A1 _21882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14935_ _24667_/Q _14933_/Y _15112_/A _24260_/Q VGND VGND VPWR VPWR _14935_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17654_ _13456_/A _16222_/C _13474_/A VGND VGND VPWR VPWR _17654_/X sky130_fd_sc_hd__o21a_4
XFILLER_36_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14866_ _14982_/A VGND VGND VPWR VPWR _14867_/A sky130_fd_sc_hd__buf_2
XFILLER_21_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22738__A _21569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16605_ _14821_/Y _16602_/X _16451_/X _16602_/X VGND VGND VPWR VPWR _16605_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21642__A _20800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13817_ _24907_/Q _24906_/Q _24905_/Q _24904_/Q VGND VGND VPWR VPWR _13817_/X sky130_fd_sc_hd__or4_4
X_17585_ _16746_/X VGND VGND VPWR VPWR _17603_/A sky130_fd_sc_hd__buf_2
XFILLER_17_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14797_ _14984_/A VGND VGND VPWR VPWR _15016_/A sky130_fd_sc_hd__buf_2
XFILLER_63_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19324_ _19323_/Y _19319_/X _19232_/X _19304_/Y VGND VGND VPWR VPWR _23375_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15640__A _15639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16536_ _16534_/Y _16530_/X _16455_/X _16535_/X VGND VGND VPWR VPWR _16536_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25041__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13748_ _24649_/Q VGND VGND VPWR VPWR _13764_/A sky130_fd_sc_hd__inv_2
XANTENNA__16538__B1 _16369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19255_ _19255_/A VGND VGND VPWR VPWR _20978_/B sky130_fd_sc_hd__inv_2
XFILLER_108_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16467_ _16467_/A VGND VGND VPWR VPWR _16467_/Y sky130_fd_sc_hd__inv_2
X_13679_ _20201_/C _13677_/X VGND VGND VPWR VPWR _13679_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__21856__A1_N _20940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18206_ _18279_/A _18278_/A _18205_/X VGND VGND VPWR VPWR _18206_/X sky130_fd_sc_hd__or3_4
X_15418_ _15418_/A _16475_/B VGND VGND VPWR VPWR _15418_/X sky130_fd_sc_hd__or2_4
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19186_ _17949_/B VGND VGND VPWR VPWR _19186_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_5_23_0_HCLK clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16398_ _16398_/A VGND VGND VPWR VPWR _16398_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22473__A _22473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18137_ _18132_/X _18137_/B _18135_/X _18136_/X VGND VGND VPWR VPWR _18164_/A sky130_fd_sc_hd__or4_4
XANTENNA__22904__C _22902_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15349_ _24605_/Q VGND VGND VPWR VPWR _22696_/A sky130_fd_sc_hd__inv_2
XFILLER_129_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22192__B _22439_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18068_ _23897_/Q VGND VGND VPWR VPWR _18068_/X sky130_fd_sc_hd__buf_2
XFILLER_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17019_ _16991_/X _17018_/X VGND VGND VPWR VPWR _17086_/A sky130_fd_sc_hd__or2_4
XFILLER_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15087__A _15087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12504__A _12403_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21598__B1 _20800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20030_ _21134_/B _20027_/X _19731_/X _20027_/X VGND VGND VPWR VPWR _20030_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15277__B1 _14236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20721__A scl_oen_o_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_147_0_HCLK clkbuf_7_73_0_HCLK/X VGND VGND VPWR VPWR _25009_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23976__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21981_ _22629_/A VGND VGND VPWR VPWR _21981_/X sky130_fd_sc_hd__buf_2
XFILLER_94_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23905__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13335__A _13334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23720_ _23753_/CLK _20530_/X HRESETn VGND VGND VPWR VPWR _23720_/Q sky130_fd_sc_hd__dfrtp_4
X_20932_ _20550_/A _11940_/Y _20741_/B _20826_/A VGND VGND VPWR VPWR _20932_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25129__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23651_ _24897_/CLK _20338_/X HRESETn VGND VGND VPWR VPWR _23651_/Q sky130_fd_sc_hd__dfrtp_4
X_20863_ _20863_/A _20863_/B _20863_/C VGND VGND VPWR VPWR _20863_/X sky130_fd_sc_hd__and3_4
XPHY_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15550__A _19448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19715__B1 _19714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22602_ _16172_/A _22524_/B VGND VGND VPWR VPWR _22602_/X sky130_fd_sc_hd__or2_4
XFILLER_126_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23582_ _23457_/CLK _23582_/D VGND VGND VPWR VPWR _17678_/B sky130_fd_sc_hd__dfxtp_4
X_20794_ _22501_/A _20787_/X _20794_/C VGND VGND VPWR VPWR _20794_/X sky130_fd_sc_hd__and3_4
XPHY_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19558__A2_N _19555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22533_ _22527_/X _22528_/X _22529_/X _22532_/X VGND VGND VPWR VPWR _22533_/X sky130_fd_sc_hd__or4_4
XFILLER_22_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13070__A _13169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22464_ _21248_/X _22463_/X _22240_/X _24517_/Q _20780_/A VGND VGND VPWR VPWR _22464_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24764__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24203_ _24244_/CLK _16442_/X HRESETn VGND VGND VPWR VPWR _16441_/A sky130_fd_sc_hd__dfrtp_4
X_21415_ _15322_/A _21414_/X _21058_/X _24505_/Q _21059_/X VGND VGND VPWR VPWR _21415_/X
+ sky130_fd_sc_hd__a32o_4
X_25183_ _25183_/CLK _11798_/X HRESETn VGND VGND VPWR VPWR _11772_/B sky130_fd_sc_hd__dfrtp_4
X_22395_ _22395_/A _22256_/B VGND VGND VPWR VPWR _22395_/X sky130_fd_sc_hd__and2_4
X_24134_ _24145_/CLK _16605_/X HRESETn VGND VGND VPWR VPWR _14821_/A sky130_fd_sc_hd__dfrtp_4
X_21346_ _21346_/A _21344_/X _21345_/X VGND VGND VPWR VPWR _21346_/X sky130_fd_sc_hd__and3_4
XANTENNA__22533__D _22532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23027__B1 _22530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21087__A2_N _20885_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12318__B2 _24493_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24065_ _24399_/CLK _16941_/X HRESETn VGND VGND VPWR VPWR _24065_/Q sky130_fd_sc_hd__dfrtp_4
X_21277_ _16121_/A _22154_/B _22351_/A VGND VGND VPWR VPWR _21277_/X sky130_fd_sc_hd__o21a_4
XFILLER_118_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23016_ _24124_/Q _22857_/B VGND VGND VPWR VPWR _23019_/B sky130_fd_sc_hd__or2_4
X_20228_ _14099_/A _20204_/X _23772_/Q VGND VGND VPWR VPWR _20264_/B sky130_fd_sc_hd__and3_4
XFILLER_46_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_43_0_HCLK clkbuf_7_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_87_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20159_ _24822_/Q _20157_/X _20158_/Y VGND VGND VPWR VPWR _20192_/B sky130_fd_sc_hd__o21a_4
XFILLER_134_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12981_ _12876_/A _12980_/X _12922_/A _12976_/B VGND VGND VPWR VPWR _12982_/A sky130_fd_sc_hd__a211o_4
XFILLER_18_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24967_ _24840_/CLK _13495_/X HRESETn VGND VGND VPWR VPWR _24967_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23646__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19954__B1 _19424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14720_ _24700_/Q VGND VGND VPWR VPWR _14876_/A sky130_fd_sc_hd__inv_2
XFILLER_45_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13245__A _13309_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11932_ _11930_/Y _11931_/X _11933_/A _11931_/X VGND VGND VPWR VPWR _25159_/D sky130_fd_sc_hd__a2bb2o_4
X_23918_ _24757_/CLK _23918_/D HRESETn VGND VGND VPWR VPWR _23918_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22558__A _21107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24898_ _24902_/CLK _13917_/X HRESETn VGND VGND VPWR VPWR _24898_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11863_ _11706_/A _11645_/X VGND VGND VPWR VPWR _11868_/A sky130_fd_sc_hd__or2_4
X_14651_ _14651_/A VGND VGND VPWR VPWR _14651_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23849_ _23845_/CLK _18325_/Y HRESETn VGND VGND VPWR VPWR _23849_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16556__A _14218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13602_ _11687_/Y _13555_/B VGND VGND VPWR VPWR _13602_/Y sky130_fd_sc_hd__nand2_4
X_17370_ _17300_/X VGND VGND VPWR VPWR _17390_/A sky130_fd_sc_hd__buf_2
XANTENNA__20316__A1 _14257_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21181__B _21638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11794_ _25184_/Q _11797_/A _11785_/X _11793_/Y VGND VGND VPWR VPWR _11794_/X sky130_fd_sc_hd__o22a_4
X_14582_ _14581_/Y VGND VGND VPWR VPWR _19144_/A sky130_fd_sc_hd__buf_2
XFILLER_25_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16321_ _16339_/A VGND VGND VPWR VPWR _16321_/X sky130_fd_sc_hd__buf_2
X_13533_ _13533_/A _13533_/B _23736_/Q _20590_/A VGND VGND VPWR VPWR _13534_/B sky130_fd_sc_hd__or4_4
XANTENNA__15397__A1_N _15395_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19040_ _13140_/B VGND VGND VPWR VPWR _19040_/Y sky130_fd_sc_hd__inv_2
X_13464_ _13403_/Y _13463_/Y _13403_/A _13463_/A VGND VGND VPWR VPWR _13464_/X sky130_fd_sc_hd__o22a_4
X_16252_ _14913_/Y _16247_/X _16251_/X _16247_/X VGND VGND VPWR VPWR _16252_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12415_ _12415_/A _12415_/B _12402_/X _12415_/D VGND VGND VPWR VPWR _12415_/X sky130_fd_sc_hd__or4_4
X_15203_ _15109_/Y _15203_/B VGND VGND VPWR VPWR _15207_/B sky130_fd_sc_hd__or2_4
XFILLER_127_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13395_ _20688_/B _13394_/X SCLK_S2 _20688_/B VGND VGND VPWR VPWR _24975_/D sky130_fd_sc_hd__a2bb2o_4
X_16183_ _16183_/A VGND VGND VPWR VPWR _16183_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24434__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16291__A _16291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12346_ _12346_/A VGND VGND VPWR VPWR _12346_/Y sky130_fd_sc_hd__inv_2
X_15134_ _15129_/A _15125_/B _15126_/X _15130_/Y VGND VGND VPWR VPWR _15135_/A sky130_fd_sc_hd__a211o_4
XANTENNA__23018__B1 _22840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18693__B1 _17199_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15065_ _15057_/X _15063_/X _15065_/C VGND VGND VPWR VPWR _24693_/D sky130_fd_sc_hd__and3_4
X_19942_ _19941_/Y _19939_/X _15561_/X _19939_/X VGND VGND VPWR VPWR _19942_/X sky130_fd_sc_hd__a2bb2o_4
X_12277_ _12176_/A _12280_/B VGND VGND VPWR VPWR _12277_/Y sky130_fd_sc_hd__nand2_4
X_14016_ _14016_/A VGND VGND VPWR VPWR _14016_/X sky130_fd_sc_hd__buf_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19873_ _23178_/Q VGND VGND VPWR VPWR _21524_/B sky130_fd_sc_hd__inv_2
X_18824_ _18821_/Y _18822_/X _18823_/X _18822_/X VGND VGND VPWR VPWR _23553_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15635__A _15431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22792__A2 _21043_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18755_ _18754_/Y _18752_/X _18685_/X _18752_/X VGND VGND VPWR VPWR _23576_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_6_0_0_HCLK clkbuf_6_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_15967_ _15965_/Y _15961_/X _11585_/X _15966_/X VGND VGND VPWR VPWR _15967_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20004__B1 _19808_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17706_ _17705_/X VGND VGND VPWR VPWR _17767_/A sky130_fd_sc_hd__inv_2
XFILLER_97_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14918_ _14918_/A _14911_/X _14918_/C _14918_/D VGND VGND VPWR VPWR _14918_/X sky130_fd_sc_hd__or4_4
XFILLER_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18686_ _18684_/Y _18682_/X _18685_/X _18682_/X VGND VGND VPWR VPWR _23600_/D sky130_fd_sc_hd__a2bb2o_4
X_15898_ _15896_/Y _15893_/X _15897_/X _15893_/X VGND VGND VPWR VPWR _15898_/X sky130_fd_sc_hd__a2bb2o_4
X_17637_ _17648_/B _17634_/Y _17636_/X _17648_/B VGND VGND VPWR VPWR _23941_/D sky130_fd_sc_hd__a2bb2o_4
X_14849_ _24688_/Q _14836_/Y _15064_/A _16601_/A VGND VGND VPWR VPWR _14849_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22187__B _22153_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24814__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17568_ _17498_/Y _17550_/B _17520_/X _17565_/Y VGND VGND VPWR VPWR _17568_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21504__B1 _21231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19307_ _23381_/Q VGND VGND VPWR VPWR _19307_/Y sky130_fd_sc_hd__inv_2
X_16519_ _16517_/Y _16518_/X _16087_/X _16518_/X VGND VGND VPWR VPWR _16519_/X sky130_fd_sc_hd__a2bb2o_4
X_17499_ _16697_/Y _17558_/B _16708_/Y _17498_/Y VGND VGND VPWR VPWR _17499_/X sky130_fd_sc_hd__or4_4
XFILLER_56_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19238_ _19238_/A VGND VGND VPWR VPWR _19238_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14537__A2 _14521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19169_ _19175_/A VGND VGND VPWR VPWR _19169_/X sky130_fd_sc_hd__buf_2
XANTENNA__24175__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14714__A _14714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21200_ _21393_/A _19005_/Y VGND VGND VPWR VPWR _21200_/X sky130_fd_sc_hd__or2_4
XANTENNA__23009__B1 _24576_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22180_ _22178_/X _22180_/B VGND VGND VPWR VPWR _22180_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__22480__B2 _16305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15529__B _15531_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24104__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22931__A _22931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15498__B1 _24560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21131_ _17629_/B VGND VGND VPWR VPWR _21348_/A sky130_fd_sc_hd__buf_2
X_21062_ _20820_/X VGND VGND VPWR VPWR _21062_/X sky130_fd_sc_hd__buf_2
XFILLER_119_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20013_ _19530_/X _19644_/X _18031_/C VGND VGND VPWR VPWR _20014_/A sky130_fd_sc_hd__or3_4
XANTENNA__18987__B2 _18982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15545__A _19445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21266__B _21043_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24821_ _23774_/CLK _14207_/X HRESETn VGND VGND VPWR VPWR _14206_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15670__B1 _11540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17760__A _14577_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21964_ _21224_/A _21960_/X _21961_/X _21962_/X _21963_/X VGND VGND VPWR VPWR _21964_/X
+ sky130_fd_sc_hd__a32o_4
X_24752_ _25009_/CLK _24752_/D HRESETn VGND VGND VPWR VPWR _14428_/A sky130_fd_sc_hd__dfstp_4
XFILLER_104_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20915_ _21860_/B _20913_/X _23036_/A _22154_/B VGND VGND VPWR VPWR _20915_/X sky130_fd_sc_hd__o22a_4
X_23703_ _23734_/CLK _20456_/Y HRESETn VGND VGND VPWR VPWR _13506_/D sky130_fd_sc_hd__dfrtp_4
XPHY_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24683_ _24712_/CLK _15093_/X HRESETn VGND VGND VPWR VPWR _24683_/Q sky130_fd_sc_hd__dfrtp_4
X_21895_ _21891_/X _21892_/X _21893_/X _21894_/X _21308_/X VGND VGND VPWR VPWR _21895_/X
+ sky130_fd_sc_hd__o41a_4
XPHY_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16376__A _16376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23634_ _23641_/CLK _23634_/D HRESETn VGND VGND VPWR VPWR _20297_/A sky130_fd_sc_hd__dfrtp_4
X_20846_ _15290_/Y _11501_/X _14096_/A _20758_/X VGND VGND VPWR VPWR _20846_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24945__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23565_ _23531_/CLK _23565_/D VGND VGND VPWR VPWR _17745_/B sky130_fd_sc_hd__dfxtp_4
X_20777_ _20749_/X VGND VGND VPWR VPWR _20777_/X sky130_fd_sc_hd__buf_2
XFILLER_11_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22516_ _22116_/X _22515_/X _21974_/X _24561_/Q _22118_/X VGND VGND VPWR VPWR _22517_/B
+ sky130_fd_sc_hd__a32o_4
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23496_ _23128_/CLK _18985_/X VGND VGND VPWR VPWR _23496_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22447_ _16520_/Y _22279_/X _24598_/Q _22170_/X VGND VGND VPWR VPWR _22447_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12200_ _25131_/Q _12200_/B VGND VGND VPWR VPWR _12200_/X sky130_fd_sc_hd__or2_4
XANTENNA__12837__A2_N _22385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13180_ _13247_/A _13176_/X _13179_/X VGND VGND VPWR VPWR _13180_/X sky130_fd_sc_hd__or3_4
X_25166_ _23898_/CLK _11876_/X HRESETn VGND VGND VPWR VPWR _11871_/A sky130_fd_sc_hd__dfrtp_4
X_22378_ _12495_/A _22259_/A _24039_/Q _22121_/X VGND VGND VPWR VPWR _22379_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_135_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15489__B1 _11563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12131_ _12123_/X _12131_/B _12131_/C _12130_/X VGND VGND VPWR VPWR _12131_/X sky130_fd_sc_hd__or4_4
XANTENNA__20482__B1 _20481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24117_ _24698_/CLK _16636_/X HRESETn VGND VGND VPWR VPWR _24117_/Q sky130_fd_sc_hd__dfrtp_4
X_21329_ _21333_/A _21329_/B VGND VGND VPWR VPWR _21330_/C sky130_fd_sc_hd__or2_4
X_25097_ _25097_/CLK _25097_/D HRESETn VGND VGND VPWR VPWR _25097_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12144__A _24573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12062_ _12062_/A VGND VGND VPWR VPWR _12062_/X sky130_fd_sc_hd__buf_2
XFILLER_2_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24048_ _24308_/CLK _24048_/D HRESETn VGND VGND VPWR VPWR _24048_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23827__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16870_ _16869_/X VGND VGND VPWR VPWR _24085_/D sky130_fd_sc_hd__inv_2
XANTENNA__16065__A1_N _16063_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15821_ _11949_/A _14195_/B _14195_/C _11514_/A VGND VGND VPWR VPWR _15821_/X sky130_fd_sc_hd__or4_4
XFILLER_65_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_130_0_HCLK clkbuf_7_65_0_HCLK/X VGND VGND VPWR VPWR _24735_/CLK sky130_fd_sc_hd__clkbuf_1
X_18540_ _18540_/A _18536_/X _18539_/Y VGND VGND VPWR VPWR _23821_/D sky130_fd_sc_hd__and3_4
XFILLER_58_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17670__A _14571_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15752_ _15757_/A VGND VGND VPWR VPWR _15752_/X sky130_fd_sc_hd__buf_2
X_12964_ _12964_/A _12964_/B VGND VGND VPWR VPWR _12964_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_193_0_HCLK clkbuf_7_96_0_HCLK/X VGND VGND VPWR VPWR _24590_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22288__A _22335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14703_ _14702_/Y VGND VGND VPWR VPWR _14703_/X sky130_fd_sc_hd__buf_2
X_11915_ _11913_/Y _11914_/X _11913_/Y _11914_/X VGND VGND VPWR VPWR _11916_/D sky130_fd_sc_hd__a2bb2o_4
X_18471_ _18470_/X VGND VGND VPWR VPWR _18472_/B sky130_fd_sc_hd__inv_2
XFILLER_46_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15683_ _12353_/Y _15680_/X _11573_/X _15680_/X VGND VGND VPWR VPWR _15683_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12895_ _12867_/X VGND VGND VPWR VPWR _12911_/A sky130_fd_sc_hd__inv_2
XFILLER_45_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17422_ _17413_/A _17413_/B VGND VGND VPWR VPWR _17422_/Y sky130_fd_sc_hd__nand2_4
X_14634_ _14633_/X _14620_/Y VGND VGND VPWR VPWR _14634_/X sky130_fd_sc_hd__and2_4
X_11846_ _19724_/A VGND VGND VPWR VPWR _19610_/A sky130_fd_sc_hd__buf_2
XANTENNA__24686__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17353_ _17353_/A _17353_/B VGND VGND VPWR VPWR _17354_/C sky130_fd_sc_hd__or2_4
XANTENNA__21920__A _21342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11777_ _11777_/A _11817_/A VGND VGND VPWR VPWR _11777_/X sky130_fd_sc_hd__and2_4
X_14565_ _14555_/X _14558_/X VGND VGND VPWR VPWR _14565_/X sky130_fd_sc_hd__and2_4
XFILLER_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24615__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16304_ _16304_/A VGND VGND VPWR VPWR _16304_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13516_ _23726_/Q _13515_/X VGND VGND VPWR VPWR _13516_/X sky130_fd_sc_hd__or2_4
X_17284_ _24006_/Q VGND VGND VPWR VPWR _17340_/A sky130_fd_sc_hd__inv_2
X_14496_ _14493_/X _14495_/X _14493_/X _14495_/X VGND VGND VPWR VPWR _14497_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA_clkbuf_4_1_0_HCLK_A clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19023_ _21505_/B _19018_/X _15559_/X _19018_/X VGND VGND VPWR VPWR _23482_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16235_ _22477_/B _16235_/B VGND VGND VPWR VPWR _16240_/A sky130_fd_sc_hd__or2_4
X_13447_ _13447_/A VGND VGND VPWR VPWR _14374_/A sky130_fd_sc_hd__inv_2
X_13378_ _13376_/Y _13372_/X _11636_/X _13377_/X VGND VGND VPWR VPWR _13378_/X sky130_fd_sc_hd__a2bb2o_4
X_16166_ _16164_/Y _16165_/X _15855_/X _16165_/X VGND VGND VPWR VPWR _24310_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15117_ _14888_/Y _14898_/Y _15117_/C VGND VGND VPWR VPWR _15117_/X sky130_fd_sc_hd__or3_4
X_12329_ _12329_/A VGND VGND VPWR VPWR _12329_/Y sky130_fd_sc_hd__inv_2
X_16097_ _16095_/Y _16090_/X _16096_/X _16090_/X VGND VGND VPWR VPWR _24336_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12054__A _12054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23006__A3 _22459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15048_ _15047_/X VGND VGND VPWR VPWR _15048_/Y sky130_fd_sc_hd__inv_2
X_19925_ _14548_/A _14543_/X _14539_/Y _19904_/D VGND VGND VPWR VPWR _19925_/X sky130_fd_sc_hd__or4_4
XFILLER_87_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15365__A _24599_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19856_ _23184_/Q VGND VGND VPWR VPWR _21215_/B sky130_fd_sc_hd__inv_2
XFILLER_84_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18807_ _18968_/A _18072_/X _18666_/C VGND VGND VPWR VPWR _18807_/X sky130_fd_sc_hd__or3_4
X_19787_ _21778_/B _19781_/X _19448_/X _19786_/X VGND VGND VPWR VPWR _23212_/D sky130_fd_sc_hd__a2bb2o_4
X_16999_ _16999_/A _16996_/X _16997_/X _16998_/X VGND VGND VPWR VPWR _16999_/X sky130_fd_sc_hd__or4_4
XANTENNA__17580__A _22395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18738_ _17750_/B VGND VGND VPWR VPWR _18738_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22198__A _22198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21725__B1 _24098_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18669_ _18664_/Y _18668_/X _17199_/X _18668_/X VGND VGND VPWR VPWR _23606_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15404__B1 _14304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20700_ _20193_/A _23616_/Q _20185_/A VGND VGND VPWR VPWR _23616_/D sky130_fd_sc_hd__a21o_4
XANTENNA__13613__A _13613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21680_ _21667_/X _19977_/Y VGND VGND VPWR VPWR _21680_/X sky130_fd_sc_hd__or2_4
X_20631_ _20630_/Y _20627_/Y VGND VGND VPWR VPWR _20631_/X sky130_fd_sc_hd__and2_4
XANTENNA__12874__D _12793_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23350_ _23350_/CLK _19398_/X VGND VGND VPWR VPWR _13030_/B sky130_fd_sc_hd__dfxtp_4
X_20562_ _20555_/A VGND VGND VPWR VPWR _20562_/X sky130_fd_sc_hd__buf_2
XFILLER_123_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20446__A _20425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22301_ _21042_/X _22300_/X _22197_/X _24406_/Q _20866_/X VGND VGND VPWR VPWR _22302_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_20_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23281_ _23303_/CLK _23281_/D VGND VGND VPWR VPWR _19587_/A sky130_fd_sc_hd__dfxtp_4
X_20493_ _20484_/X _20492_/X _15363_/A _20488_/X VGND VGND VPWR VPWR _23711_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25020_ _25021_/CLK _12959_/X HRESETn VGND VGND VPWR VPWR _22474_/A sky130_fd_sc_hd__dfrtp_4
X_22232_ _22232_/A _22265_/B VGND VGND VPWR VPWR _22232_/X sky130_fd_sc_hd__and2_4
XANTENNA__17238__A2_N _25221_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22083__D _22082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22453__B2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14930__A2 _24273_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12941__A1 _12854_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22163_ _22163_/A _22160_/X _22162_/X VGND VGND VPWR VPWR _22163_/X sky130_fd_sc_hd__and3_4
XFILLER_117_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16132__A1 _15421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23991__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21114_ _21113_/X VGND VGND VPWR VPWR _21867_/A sky130_fd_sc_hd__buf_2
X_22094_ _22087_/A _22094_/B VGND VGND VPWR VPWR _22094_/X sky130_fd_sc_hd__or2_4
XFILLER_120_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23920__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15891__B1 _15890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21045_ _21034_/Y VGND VGND VPWR VPWR _22197_/A sky130_fd_sc_hd__buf_2
XFILLER_99_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19082__B1 _19038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25144__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13507__B _13506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22508__A2 _22574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17490__A _17490_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24804_ _24811_/CLK _14256_/X HRESETn VGND VGND VPWR VPWR _14255_/A sky130_fd_sc_hd__dfstp_4
Xclkbuf_8_203_0_HCLK clkbuf_8_203_0_HCLK/A VGND VGND VPWR VPWR _24055_/CLK sky130_fd_sc_hd__clkbuf_1
X_22996_ _22995_/X VGND VGND VPWR VPWR _22996_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_9_0_HCLK clkbuf_7_4_0_HCLK/X VGND VGND VPWR VPWR _23939_/CLK sky130_fd_sc_hd__clkbuf_1
X_24735_ _24735_/CLK _24735_/D HRESETn VGND VGND VPWR VPWR _17717_/A sky130_fd_sc_hd__dfrtp_4
X_21947_ _21393_/A _21947_/B VGND VGND VPWR VPWR _21947_/X sky130_fd_sc_hd__or2_4
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17396__B1 _17345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11700_ _11698_/D VGND VGND VPWR VPWR _18638_/B sky130_fd_sc_hd__inv_2
XPHY_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12679_/X VGND VGND VPWR VPWR _12685_/B sky130_fd_sc_hd__inv_2
XPHY_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21878_ _13630_/C _21875_/X _21877_/X VGND VGND VPWR VPWR _21878_/X sky130_fd_sc_hd__and3_4
XPHY_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24666_ _24671_/CLK _15180_/X HRESETn VGND VGND VPWR VPWR _14894_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _15282_/A VGND VGND VPWR VPWR _11631_/X sky130_fd_sc_hd__buf_2
XFILLER_42_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ _21591_/B VGND VGND VPWR VPWR _22859_/A sky130_fd_sc_hd__buf_2
XPHY_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23617_ _24783_/CLK _23617_/D HRESETn VGND VGND VPWR VPWR _23617_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23774__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24097__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22141__B1 _21581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24597_ _24055_/CLK _15372_/X HRESETn VGND VGND VPWR VPWR _15371_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11562_ _11562_/A VGND VGND VPWR VPWR _11562_/Y sky130_fd_sc_hd__inv_2
X_14350_ _13845_/X VGND VGND VPWR VPWR _14350_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23548_ _23482_/CLK _23548_/D VGND VGND VPWR VPWR _23548_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13301_ _13301_/A _23199_/Q VGND VGND VPWR VPWR _13302_/C sky130_fd_sc_hd__or2_4
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14281_ _14279_/Y _14280_/X _14213_/X _14280_/X VGND VGND VPWR VPWR _14281_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11978__A _11965_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23479_ _23479_/CLK _23479_/D VGND VGND VPWR VPWR _19029_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13232_ _13232_/A _13228_/X _13231_/X VGND VGND VPWR VPWR _13232_/X sky130_fd_sc_hd__or3_4
X_16020_ _16016_/X VGND VGND VPWR VPWR _16020_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21247__A2 _21244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25218_ _24405_/CLK _11538_/X HRESETn VGND VGND VPWR VPWR _25218_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20455__B1 _20446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13163_ _13159_/X _13161_/X _13162_/X VGND VGND VPWR VPWR _13164_/C sky130_fd_sc_hd__and3_4
X_25149_ _24851_/CLK _25149_/D HRESETn VGND VGND VPWR VPWR _11980_/A sky130_fd_sc_hd__dfrtp_4
X_12114_ _24547_/Q VGND VGND VPWR VPWR _12114_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21187__A _22198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13094_ _13137_/A _23365_/Q VGND VGND VPWR VPWR _13094_/X sky130_fd_sc_hd__or2_4
X_17971_ _15729_/X _17955_/X _17970_/X _23927_/Q _15728_/A VGND VGND VPWR VPWR _17971_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__23661__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19710_ _19709_/Y VGND VGND VPWR VPWR _19710_/X sky130_fd_sc_hd__buf_2
X_12045_ _12045_/A _12045_/B _12045_/C _12044_/X VGND VGND VPWR VPWR _12045_/X sky130_fd_sc_hd__or4_4
X_16922_ _16922_/A _16922_/B VGND VGND VPWR VPWR _16942_/A sky130_fd_sc_hd__or2_4
XFILLER_46_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_13_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19641_ _25169_/Q VGND VGND VPWR VPWR _19641_/X sky130_fd_sc_hd__buf_2
XFILLER_78_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16853_ _16853_/A _16853_/B VGND VGND VPWR VPWR _16854_/A sky130_fd_sc_hd__or2_4
XANTENNA__21915__A _21930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18820__B1 _18795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15634__B1 _14304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15804_ _15799_/X _15582_/A _15735_/X _20834_/A _15746_/A VGND VGND VPWR VPWR _24429_/D
+ sky130_fd_sc_hd__a32o_4
X_19572_ _19571_/Y _19567_/X _19256_/X _19554_/Y VGND VGND VPWR VPWR _19572_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15913__A _15916_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16784_ _16784_/A VGND VGND VPWR VPWR _16784_/Y sky130_fd_sc_hd__inv_2
X_13996_ _24810_/Q VGND VGND VPWR VPWR _13996_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18523_ _18485_/C _18427_/C VGND VGND VPWR VPWR _18523_/X sky130_fd_sc_hd__or2_4
X_15735_ _15431_/X VGND VGND VPWR VPWR _15735_/X sky130_fd_sc_hd__buf_2
XFILLER_20_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12947_ _12947_/A _12947_/B VGND VGND VPWR VPWR _12947_/X sky130_fd_sc_hd__or2_4
XFILLER_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21183__B2 _21716_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18454_ _23842_/Q _18453_/Y VGND VGND VPWR VPWR _18454_/X sky130_fd_sc_hd__or2_4
XFILLER_45_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15666_ _15666_/A VGND VGND VPWR VPWR _15666_/X sky130_fd_sc_hd__buf_2
XFILLER_60_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12878_ _12878_/A _12878_/B _12878_/C _12974_/A VGND VGND VPWR VPWR _12933_/D sky130_fd_sc_hd__or4_4
XANTENNA__20930__A1 _20910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14248__B _18633_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17405_ _17325_/B _17399_/X _17401_/Y _17336_/X VGND VGND VPWR VPWR _17406_/A sky130_fd_sc_hd__a211o_4
X_14617_ _14608_/Y _14615_/Y _14617_/C VGND VGND VPWR VPWR _14617_/X sky130_fd_sc_hd__and3_4
X_11829_ _11815_/C _11809_/B _11828_/X VGND VGND VPWR VPWR _11830_/A sky130_fd_sc_hd__or3_4
X_18385_ _16438_/Y _23827_/Q _16438_/Y _23827_/Q VGND VGND VPWR VPWR _18385_/X sky130_fd_sc_hd__a2bb2o_4
X_15597_ _15574_/X _15582_/X _15596_/X _24527_/Q _15585_/X VGND VGND VPWR VPWR _15597_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_18_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _17622_/B VGND VGND VPWR VPWR _17336_/X sky130_fd_sc_hd__buf_2
XANTENNA__19120__A _18711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14548_ _14548_/A VGND VGND VPWR VPWR _14548_/X sky130_fd_sc_hd__buf_2
XFILLER_81_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18887__B1 _18817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22683__B2 _22322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17267_ _11568_/A _23996_/Q _11568_/Y _17266_/Y VGND VGND VPWR VPWR _17267_/X sky130_fd_sc_hd__o22a_4
XFILLER_35_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14479_ _14479_/A VGND VGND VPWR VPWR _14480_/A sky130_fd_sc_hd__inv_2
XFILLER_128_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19006_ _19005_/Y _19003_/X _15566_/X _19003_/X VGND VGND VPWR VPWR _23488_/D sky130_fd_sc_hd__a2bb2o_4
X_16218_ _24289_/Q VGND VGND VPWR VPWR _16218_/Y sky130_fd_sc_hd__inv_2
X_17198_ _17213_/A VGND VGND VPWR VPWR _17198_/X sky130_fd_sc_hd__buf_2
XFILLER_122_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23749__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16149_ _24316_/Q VGND VGND VPWR VPWR _16149_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22199__B1 _24404_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15095__A _15158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19908_ _19908_/A VGND VGND VPWR VPWR _21962_/B sky130_fd_sc_hd__inv_2
XFILLER_114_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21825__A _20975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19839_ _19839_/A VGND VGND VPWR VPWR _22057_/B sky130_fd_sc_hd__inv_2
XFILLER_111_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13327__B _21707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15625__B1 _15513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22850_ _21546_/X _22846_/Y _22423_/X _22849_/X VGND VGND VPWR VPWR _22851_/D sky130_fd_sc_hd__a2bb2o_4
X_21801_ _21801_/A _20072_/Y _21800_/X VGND VGND VPWR VPWR _21801_/X sky130_fd_sc_hd__and3_4
X_22781_ _22418_/X _22781_/B _22781_/C VGND VGND VPWR VPWR _22781_/X sky130_fd_sc_hd__and3_4
XANTENNA__17378__B1 _17345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24537__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22371__B1 _24407_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21732_ _21731_/X VGND VGND VPWR VPWR _21732_/Y sky130_fd_sc_hd__inv_2
X_24520_ _24521_/CLK _15609_/X HRESETn VGND VGND VPWR VPWR _12588_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_33_0_HCLK clkbuf_8_33_0_HCLK/A VGND VGND VPWR VPWR _23288_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__11662__B2 _23917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_96_0_HCLK clkbuf_7_48_0_HCLK/X VGND VGND VPWR VPWR _24071_/CLK sky130_fd_sc_hd__clkbuf_1
X_21663_ _21657_/A _21663_/B VGND VGND VPWR VPWR _21663_/X sky130_fd_sc_hd__or2_4
XFILLER_75_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24451_ _24451_/CLK _24451_/D HRESETn VGND VGND VPWR VPWR _12853_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24190__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20614_ _13535_/X VGND VGND VPWR VPWR _20614_/Y sky130_fd_sc_hd__inv_2
X_23402_ _23112_/CLK _23402_/D VGND VGND VPWR VPWR _23402_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18878__B1 _18764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24382_ _24378_/CLK _24382_/D HRESETn VGND VGND VPWR VPWR _24382_/Q sky130_fd_sc_hd__dfrtp_4
X_21594_ _17027_/A _13333_/A VGND VGND VPWR VPWR _21594_/X sky130_fd_sc_hd__or2_4
XFILLER_36_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23333_ _23313_/CLK _19446_/X VGND VGND VPWR VPWR _23333_/Q sky130_fd_sc_hd__dfxtp_4
X_20545_ _20545_/A VGND VGND VPWR VPWR _20545_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22426__A1 _24559_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23264_ _23249_/CLK _23264_/D VGND VGND VPWR VPWR _23264_/Q sky130_fd_sc_hd__dfxtp_4
X_20476_ _20461_/X _20475_/X _15373_/A _20466_/X VGND VGND VPWR VPWR _23707_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22391__A _24480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22215_ _22215_/A _12065_/A VGND VGND VPWR VPWR _22215_/Y sky130_fd_sc_hd__nor2_4
X_25003_ _25002_/CLK _13056_/X HRESETn VGND VGND VPWR VPWR _25003_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17485__A _22307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23195_ _23154_/CLK _23195_/D VGND VGND VPWR VPWR _23195_/Q sky130_fd_sc_hd__dfxtp_4
X_22146_ _14726_/A _22146_/B VGND VGND VPWR VPWR _22146_/X sky130_fd_sc_hd__or2_4
XFILLER_117_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22077_ _21764_/A _22075_/X _22076_/X VGND VGND VPWR VPWR _22077_/X sky130_fd_sc_hd__and3_4
XANTENNA__12422__A _12434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21028_ _20772_/Y _21028_/B _20898_/Y _21027_/Y VGND VGND VPWR VPWR HRDATA[0] sky130_fd_sc_hd__or4_4
XFILLER_43_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15616__B1 _24515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13850_ _13815_/X _13812_/X VGND VGND VPWR VPWR _13872_/C sky130_fd_sc_hd__or2_4
XFILLER_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24960__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12801_ _22160_/A _22161_/A _12984_/A _12800_/Y VGND VGND VPWR VPWR _12801_/X sky130_fd_sc_hd__o22a_4
X_13781_ _13726_/X _13728_/X _13730_/X _13732_/D VGND VGND VPWR VPWR _13781_/X sky130_fd_sc_hd__or4_4
XANTENNA__24278__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22362__B1 _25202_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22979_ _22979_/A _23004_/A VGND VGND VPWR VPWR _22982_/B sky130_fd_sc_hd__and2_4
X_15520_ _11625_/A VGND VGND VPWR VPWR _15520_/X sky130_fd_sc_hd__buf_2
X_12732_ _12749_/A _12732_/B _12732_/C VGND VGND VPWR VPWR _25050_/D sky130_fd_sc_hd__and3_4
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18046__A1_N _21335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24718_ _23664_/CLK _24718_/D HRESETn VGND VGND VPWR VPWR _24718_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20018__A2_N _20015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24207__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21470__A _21336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15451_ _14432_/A _15453_/A _15443_/X _15450_/Y VGND VGND VPWR VPWR _24578_/D sky130_fd_sc_hd__o22a_4
XFILLER_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12663_ _12663_/A _12663_/B VGND VGND VPWR VPWR _12663_/X sky130_fd_sc_hd__or2_4
XFILLER_15_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24649_ _24641_/CLK _24649_/D HRESETn VGND VGND VPWR VPWR _24649_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16564__A _23008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _13432_/Y _14402_/B VGND VGND VPWR VPWR _14402_/Y sky130_fd_sc_hd__nand2_4
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _11614_/A VGND VGND VPWR VPWR _11614_/Y sky130_fd_sc_hd__inv_2
X_18170_ _16095_/Y _18209_/A _16095_/Y _18209_/A VGND VGND VPWR VPWR _18172_/C sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_5_4_0_HCLK clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15382_ _22212_/A _15381_/X _11604_/X _15381_/X VGND VGND VPWR VPWR _24593_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22716__D _22715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _25054_/Q _12592_/Y _12593_/Y _12596_/A VGND VGND VPWR VPWR _12594_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17121_ _17116_/A _17116_/B _17083_/X _17117_/Y VGND VGND VPWR VPWR _17122_/A sky130_fd_sc_hd__a211o_4
XFILLER_51_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14333_ _24778_/Q _14325_/X _24777_/Q _14327_/X VGND VGND VPWR VPWR _14333_/X sky130_fd_sc_hd__o22a_4
X_11545_ HWDATA[26] VGND VGND VPWR VPWR _11545_/X sky130_fd_sc_hd__buf_2
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17052_ _17052_/A _17050_/X _17051_/Y VGND VGND VPWR VPWR _24058_/D sky130_fd_sc_hd__and3_4
X_14264_ _24800_/Q VGND VGND VPWR VPWR _14264_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16003_ _15435_/A VGND VGND VPWR VPWR _16003_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23842__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13215_ _13247_/A _13211_/X _13214_/X VGND VGND VPWR VPWR _13215_/X sky130_fd_sc_hd__or3_4
XFILLER_124_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25066__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14195_ _11949_/A _14195_/B _14195_/C _16038_/D VGND VGND VPWR VPWR _21072_/A sky130_fd_sc_hd__or4_4
XFILLER_83_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13146_ _13146_/A _13146_/B VGND VGND VPWR VPWR _13147_/C sky130_fd_sc_hd__or2_4
XFILLER_124_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17240__A1_N _11614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13428__A _13428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13077_ _13127_/A _23075_/Q VGND VGND VPWR VPWR _13080_/B sky130_fd_sc_hd__or2_4
X_17954_ _17725_/A _17954_/B _17954_/C VGND VGND VPWR VPWR _17955_/C sky130_fd_sc_hd__or3_4
X_12028_ _11999_/A _12027_/Y _11999_/A _12027_/Y VGND VGND VPWR VPWR _12028_/X sky130_fd_sc_hd__a2bb2o_4
X_16905_ _16890_/A _16902_/B _16904_/Y VGND VGND VPWR VPWR _24075_/D sky130_fd_sc_hd__and3_4
X_17885_ _17853_/A _19181_/A VGND VGND VPWR VPWR _17886_/C sky130_fd_sc_hd__or2_4
XFILLER_120_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15643__A _15642_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16836_ _24059_/Q VGND VGND VPWR VPWR _16837_/D sky130_fd_sc_hd__inv_2
X_19624_ _19636_/A VGND VGND VPWR VPWR _19624_/X sky130_fd_sc_hd__buf_2
XANTENNA__19115__A _11635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16280__B1 _16279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19555_ _19554_/Y VGND VGND VPWR VPWR _19555_/X sky130_fd_sc_hd__buf_2
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16767_ _24067_/Q VGND VGND VPWR VPWR _16935_/A sky130_fd_sc_hd__inv_2
X_13979_ _13971_/X _13978_/Y _24888_/Q _13971_/X VGND VGND VPWR VPWR _13979_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22353__B1 _20799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18506_ _18506_/A VGND VGND VPWR VPWR _23829_/D sky130_fd_sc_hd__inv_2
X_15718_ _15717_/X VGND VGND VPWR VPWR _15718_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19486_ _23318_/Q VGND VGND VPWR VPWR _19486_/Y sky130_fd_sc_hd__inv_2
X_16698_ _22598_/A _23960_/Q _15955_/Y _16697_/Y VGND VGND VPWR VPWR _16698_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12841__B1 _22712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22476__A _21246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18437_ _18469_/A _18468_/A _18437_/C _18468_/B VGND VGND VPWR VPWR _18438_/B sky130_fd_sc_hd__or4_4
X_15649_ _15411_/X _15647_/X _15635_/X _24500_/Q _15648_/X VGND VGND VPWR VPWR _24500_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_61_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18368_ _23832_/Q VGND VGND VPWR VPWR _18434_/C sky130_fd_sc_hd__inv_2
X_17319_ _17319_/A VGND VGND VPWR VPWR _17319_/Y sky130_fd_sc_hd__inv_2
X_18299_ _16296_/Y _18299_/B VGND VGND VPWR VPWR _18299_/X sky130_fd_sc_hd__or2_4
XFILLER_119_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22923__B _22920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20330_ _14266_/X _20330_/B VGND VGND VPWR VPWR _20330_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__14346__B1 _23077_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12606__A2_N _24525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20261_ _20212_/D VGND VGND VPWR VPWR _20264_/A sky130_fd_sc_hd__inv_2
XFILLER_134_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14722__A _14722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22000_ _15456_/X VGND VGND VPWR VPWR _22259_/A sky130_fd_sc_hd__buf_2
XFILLER_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20192_ _20192_/A _20192_/B VGND VGND VPWR VPWR _20192_/X sky130_fd_sc_hd__and2_4
XFILLER_88_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13338__A _14047_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24789__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13321__B2 _13054_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23951_ _24079_/CLK _17601_/X HRESETn VGND VGND VPWR VPWR _22202_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24718__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22592__B1 _12117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15553__A _19455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22902_ _16693_/A _22654_/X _22564_/B VGND VGND VPWR VPWR _22902_/X sky130_fd_sc_hd__a21o_4
XANTENNA__21274__B _22444_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23882_ _23885_/CLK _23882_/D HRESETn VGND VGND VPWR VPWR _18120_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_56_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_4_0_HCLK_A clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16271__B1 _24271_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15613__A3 _15494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22833_ _22249_/A VGND VGND VPWR VPWR _22834_/B sky130_fd_sc_hd__buf_2
XFILLER_38_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24371__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13073__A _13073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22895__A1 _21572_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24300__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22764_ _21572_/B _22763_/X _22640_/X _25213_/Q _22641_/X VGND VGND VPWR VPWR _22764_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24503_ _25009_/CLK _15634_/X HRESETn VGND VGND VPWR VPWR _24503_/Q sky130_fd_sc_hd__dfrtp_4
X_21715_ _16300_/A VGND VGND VPWR VPWR _21715_/X sky130_fd_sc_hd__buf_2
XFILLER_24_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16574__A1 _15799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22695_ _22695_/A _22435_/X VGND VGND VPWR VPWR _22695_/X sky130_fd_sc_hd__and2_4
XFILLER_129_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21646_ _21643_/X _21644_/X _21645_/X VGND VGND VPWR VPWR _21646_/Y sky130_fd_sc_hd__o21ai_4
X_24434_ _25012_/CLK _24434_/D HRESETn VGND VGND VPWR VPWR _21851_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_36_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20658__B1 _20583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21577_ _21575_/Y _21576_/X _13503_/A _21020_/B VGND VGND VPWR VPWR _21577_/X sky130_fd_sc_hd__a2bb2o_4
X_24365_ _24405_/CLK _24365_/D HRESETn VGND VGND VPWR VPWR _24365_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12417__A _12417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20528_ _23720_/Q _20524_/A _20524_/B VGND VGND VPWR VPWR _20528_/X sky130_fd_sc_hd__or3_4
X_23316_ _23313_/CLK _19495_/X VGND VGND VPWR VPWR _19493_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_125_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24296_ _24031_/CLK _24296_/D HRESETn VGND VGND VPWR VPWR _16200_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18079__A1 _21188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20459_ _22212_/A _20437_/X _20446_/X _20458_/X VGND VGND VPWR VPWR _20460_/A sky130_fd_sc_hd__o22a_4
XFILLER_4_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23247_ _23356_/CLK _19685_/X VGND VGND VPWR VPWR _19684_/A sky130_fd_sc_hd__dfxtp_4
X_13000_ _12818_/Y _12999_/X VGND VGND VPWR VPWR _13004_/B sky130_fd_sc_hd__or2_4
XFILLER_107_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23178_ _23156_/CLK _23178_/D VGND VGND VPWR VPWR _23178_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11571__B1 _11570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22129_ _20783_/X VGND VGND VPWR VPWR _22129_/X sky130_fd_sc_hd__buf_2
XANTENNA__13248__A _13092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17943__A _17732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12115__A2 _24547_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14951_ _14950_/Y _22477_/A _14950_/Y _22477_/A VGND VGND VPWR VPWR _14951_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16559__A _16559_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24459__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13902_ _13824_/X _13892_/X _13884_/X _13867_/A _13893_/X VGND VGND VPWR VPWR _24908_/D
+ sky130_fd_sc_hd__a32o_4
X_17670_ _14571_/X VGND VGND VPWR VPWR _17697_/A sky130_fd_sc_hd__buf_2
X_14882_ _14882_/A _14881_/X VGND VGND VPWR VPWR _14987_/A sky130_fd_sc_hd__or2_4
XFILLER_63_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16621_ _16621_/A _16235_/B VGND VGND VPWR VPWR _16627_/A sky130_fd_sc_hd__or2_4
X_13833_ _13833_/A _13869_/B _24904_/Q _13833_/D VGND VGND VPWR VPWR _13833_/X sky130_fd_sc_hd__and4_4
XFILLER_1_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19340_ _13241_/B VGND VGND VPWR VPWR _19340_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16552_ _16551_/Y _16549_/X _16291_/X _16549_/X VGND VGND VPWR VPWR _24160_/D sky130_fd_sc_hd__a2bb2o_4
X_13764_ _13764_/A VGND VGND VPWR VPWR _13764_/X sky130_fd_sc_hd__buf_2
XANTENNA__24041__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15503_ _11532_/X VGND VGND VPWR VPWR _15503_/X sky130_fd_sc_hd__buf_2
XFILLER_95_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12715_ _12587_/Y _12714_/X VGND VGND VPWR VPWR _12715_/Y sky130_fd_sc_hd__nand2_4
X_19271_ _21756_/B VGND VGND VPWR VPWR _19271_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19751__B2 _19750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16483_ _24187_/Q VGND VGND VPWR VPWR _16483_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15910__B _16127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13695_ _24920_/Q _13687_/X _21733_/A _13689_/X VGND VGND VPWR VPWR _13695_/X sky130_fd_sc_hd__o22a_4
X_18222_ _18258_/A _18222_/B _18179_/Y _18222_/D VGND VGND VPWR VPWR _18223_/B sky130_fd_sc_hd__or4_4
XFILLER_31_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15434_ _15430_/X _15415_/Y _15432_/X _13546_/A _15433_/X VGND VGND VPWR VPWR _15434_/X
+ sky130_fd_sc_hd__a32o_4
X_12646_ _12704_/A _12701_/A _12700_/A VGND VGND VPWR VPWR _12646_/X sky130_fd_sc_hd__or3_4
XFILLER_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18153_ _24331_/Q _18152_/A _22014_/A _18316_/A VGND VGND VPWR VPWR _18153_/X sky130_fd_sc_hd__o22a_4
X_15365_ _24599_/Q VGND VGND VPWR VPWR _22487_/A sky130_fd_sc_hd__inv_2
X_12577_ _12577_/A _12570_/X _12577_/C _12576_/X VGND VGND VPWR VPWR _12591_/C sky130_fd_sc_hd__or4_4
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21310__B2 _21113_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17104_ _17042_/A _16992_/Y _17042_/D _17096_/B VGND VGND VPWR VPWR _17104_/X sky130_fd_sc_hd__or4_4
XFILLER_117_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14316_ _23649_/Q VGND VGND VPWR VPWR _14329_/A sky130_fd_sc_hd__buf_2
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ _11527_/Y VGND VGND VPWR VPWR _11529_/A sky130_fd_sc_hd__buf_2
X_18084_ _11749_/X _18086_/A _18081_/X VGND VGND VPWR VPWR _18084_/X sky130_fd_sc_hd__o21a_4
X_15296_ HTRANS[1] VGND VGND VPWR VPWR _15296_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17007__A2_N _17027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17035_ _17133_/A _17029_/X _17035_/C _17034_/X VGND VGND VPWR VPWR _17124_/B sky130_fd_sc_hd__or4_4
X_14247_ _14247_/A VGND VGND VPWR VPWR _14247_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15638__A _15637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19267__B1 _19152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21074__B1 _24801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14178_ _14175_/X _14177_/Y _25155_/Q _14175_/X VGND VGND VPWR VPWR _24831_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13129_ _13203_/A _13129_/B _13128_/X VGND VGND VPWR VPWR _13133_/B sky130_fd_sc_hd__and3_4
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18986_ _18986_/A VGND VGND VPWR VPWR _18986_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24882__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17937_ _17969_/A _17937_/B _17936_/X VGND VGND VPWR VPWR _17937_/X sky130_fd_sc_hd__or3_4
XFILLER_61_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17868_ _17796_/X _17868_/B VGND VGND VPWR VPWR _17869_/C sky130_fd_sc_hd__or2_4
XANTENNA__24129__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16253__B1 _24278_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19607_ _19607_/A VGND VGND VPWR VPWR _19607_/X sky130_fd_sc_hd__buf_2
XFILLER_53_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16819_ _24085_/Q VGND VGND VPWR VPWR _16819_/Y sky130_fd_sc_hd__inv_2
X_17799_ _14571_/X _18926_/A VGND VGND VPWR VPWR _17799_/X sky130_fd_sc_hd__or2_4
XFILLER_93_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19538_ _23300_/Q VGND VGND VPWR VPWR _19538_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11908__A1_N _11904_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20888__B1 _12011_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19469_ _19466_/Y _19468_/X _17993_/X _19468_/X VGND VGND VPWR VPWR _19469_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21500_ _21500_/A _21498_/X _21499_/X VGND VGND VPWR VPWR _21500_/X sky130_fd_sc_hd__and3_4
X_22480_ _22264_/X _22479_/X _16349_/Y _16305_/X VGND VGND VPWR VPWR _22480_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14436__B _14436_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23764__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21431_ _24292_/Q _21293_/B VGND VGND VPWR VPWR _21431_/X sky130_fd_sc_hd__or2_4
XFILLER_124_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_107_0_HCLK clkbuf_7_53_0_HCLK/X VGND VGND VPWR VPWR _24620_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12545__A2_N _24533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21301__A1 _14818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16932__A _16936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24150_ _24104_/CLK _24150_/D HRESETn VGND VGND VPWR VPWR _24150_/Q sky130_fd_sc_hd__dfrtp_4
X_21362_ _21357_/X _21361_/X _11688_/Y _21357_/X VGND VGND VPWR VPWR _21362_/X sky130_fd_sc_hd__a2bb2o_4
X_20313_ _20313_/A VGND VGND VPWR VPWR _20313_/Y sky130_fd_sc_hd__inv_2
X_23101_ _23278_/CLK _20078_/X VGND VGND VPWR VPWR _20074_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__19773__A2_N _19772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24081_ _24064_/CLK _16882_/Y HRESETn VGND VGND VPWR VPWR _24081_/Q sky130_fd_sc_hd__dfrtp_4
X_21293_ _21293_/A _21293_/B VGND VGND VPWR VPWR _21293_/X sky130_fd_sc_hd__or2_4
X_23032_ _14366_/X _23032_/B VGND VGND VPWR VPWR _23759_/D sky130_fd_sc_hd__or2_4
X_20244_ _20244_/A _20225_/B VGND VGND VPWR VPWR _20244_/X sky130_fd_sc_hd__and2_4
XFILLER_116_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11553__B1 _11552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17763__A _16678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20175_ _20175_/A VGND VGND VPWR VPWR _20234_/B sky130_fd_sc_hd__buf_2
XFILLER_27_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24552__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24983_ _24984_/CLK _24983_/D HRESETn VGND VGND VPWR VPWR _13368_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_130_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23934_ _23486_/CLK _17669_/X HRESETn VGND VGND VPWR VPWR _13406_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_57_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16244__B1 _16243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23865_ _23859_/CLK _18271_/Y HRESETn VGND VGND VPWR VPWR _23865_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_38_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17992__B1 _16455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22816_ _22681_/A _22816_/B VGND VGND VPWR VPWR _22816_/X sky130_fd_sc_hd__and2_4
XANTENNA__22868__B2 _22531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23796_ _23796_/CLK _23796_/D HRESETn VGND VGND VPWR VPWR _23796_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23005__A _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22747_ _24148_/Q _22505_/X _22576_/X _22746_/X VGND VGND VPWR VPWR _22748_/C sky130_fd_sc_hd__a211o_4
XFILLER_73_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12500_ _12495_/A _12495_/B _12453_/X _12497_/B VGND VGND VPWR VPWR _12500_/X sky130_fd_sc_hd__a211o_4
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13480_ _13480_/A _13480_/B VGND VGND VPWR VPWR _13480_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_66_0_HCLK clkbuf_7_67_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_66_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22678_ _22678_/A _22956_/B VGND VGND VPWR VPWR _22681_/B sky130_fd_sc_hd__or2_4
XFILLER_40_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22844__A _24455_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12431_ _12433_/B VGND VGND VPWR VPWR _12432_/B sky130_fd_sc_hd__inv_2
X_24417_ _24425_/CLK _24417_/D HRESETn VGND VGND VPWR VPWR _24417_/Q sky130_fd_sc_hd__dfrtp_4
X_21629_ _21617_/A _21629_/B VGND VGND VPWR VPWR _21629_/X sky130_fd_sc_hd__or2_4
XFILLER_138_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15150_ _15138_/B _15154_/B VGND VGND VPWR VPWR _15151_/C sky130_fd_sc_hd__nand2_4
X_12362_ _12362_/A VGND VGND VPWR VPWR _12411_/B sky130_fd_sc_hd__inv_2
X_24348_ _24333_/CLK _24348_/D HRESETn VGND VGND VPWR VPWR _16063_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14101_ _23770_/Q VGND VGND VPWR VPWR _20200_/A sky130_fd_sc_hd__buf_2
X_12293_ _12265_/A _12293_/B VGND VGND VPWR VPWR _12293_/Y sky130_fd_sc_hd__nand2_4
X_15081_ _24687_/Q _15080_/Y VGND VGND VPWR VPWR _15081_/X sky130_fd_sc_hd__or2_4
X_24279_ _24681_/CLK _16252_/X HRESETn VGND VGND VPWR VPWR _24279_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12336__A2 _24474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14032_ _20209_/A VGND VGND VPWR VPWR _20246_/A sky130_fd_sc_hd__inv_2
XFILLER_122_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17673__A _14569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18840_ _23547_/Q VGND VGND VPWR VPWR _18840_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18771_ _18771_/A VGND VGND VPWR VPWR _18771_/Y sky130_fd_sc_hd__inv_2
X_15983_ _15981_/Y _15979_/X _15982_/X _15979_/X VGND VGND VPWR VPWR _24368_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24293__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17722_ _17881_/A _23149_/Q VGND VGND VPWR VPWR _17723_/C sky130_fd_sc_hd__or2_4
X_14934_ _15218_/A VGND VGND VPWR VPWR _15112_/A sky130_fd_sc_hd__inv_2
XFILLER_76_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24222__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17432__C1 _17345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17653_ _13407_/A VGND VGND VPWR VPWR _17653_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21923__A _17636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14865_ _14864_/X VGND VGND VPWR VPWR _14865_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16604_ _14831_/Y _16602_/X _16279_/X _16602_/X VGND VGND VPWR VPWR _16604_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13816_ _13816_/A VGND VGND VPWR VPWR _13867_/A sky130_fd_sc_hd__buf_2
X_17584_ _17583_/X VGND VGND VPWR VPWR _17584_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16250__A3 _15596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14796_ _14982_/A VGND VGND VPWR VPWR _14984_/A sky130_fd_sc_hd__inv_2
X_19323_ _13309_/B VGND VGND VPWR VPWR _19323_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16535_ _16530_/A VGND VGND VPWR VPWR _16535_/X sky130_fd_sc_hd__buf_2
X_13747_ _13716_/B VGND VGND VPWR VPWR _13769_/B sky130_fd_sc_hd__buf_2
X_19254_ _21169_/B _19251_/X _11860_/X _19251_/X VGND VGND VPWR VPWR _23400_/D sky130_fd_sc_hd__a2bb2o_4
X_16466_ _16464_/Y _16460_/X _15992_/X _16465_/X VGND VGND VPWR VPWR _24194_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13678_ _23687_/Q VGND VGND VPWR VPWR _13678_/X sky130_fd_sc_hd__buf_2
X_18205_ _18205_/A _18202_/Y _18203_/Y _18205_/D VGND VGND VPWR VPWR _18205_/X sky130_fd_sc_hd__or4_4
X_15417_ _14197_/A VGND VGND VPWR VPWR _15418_/A sky130_fd_sc_hd__buf_2
X_12629_ _12629_/A VGND VGND VPWR VPWR _12629_/X sky130_fd_sc_hd__buf_2
X_19185_ _19184_/Y _19182_/X _19095_/X _19182_/X VGND VGND VPWR VPWR _23424_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25081__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16397_ _16389_/Y _16396_/X _15320_/X _16396_/X VGND VGND VPWR VPWR _16397_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18136_ _16061_/Y _18199_/A _16061_/Y _18199_/A VGND VGND VPWR VPWR _18136_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21295__B1 _20744_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15348_ _15347_/Y _15345_/X _11558_/X _15345_/X VGND VGND VPWR VPWR _15348_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25010__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22904__D _22903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18067_ _18067_/A VGND VGND VPWR VPWR _18067_/X sky130_fd_sc_hd__buf_2
XFILLER_32_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15368__A _11532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15279_ _13632_/A VGND VGND VPWR VPWR _15279_/X sky130_fd_sc_hd__buf_2
XFILLER_67_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17018_ _16999_/X _17004_/X _17012_/X _17017_/X VGND VGND VPWR VPWR _17018_/X sky130_fd_sc_hd__or4_4
XFILLER_125_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21598__A1 _21064_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22795__B1 _16157_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18679__A _18678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24837__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13319__C _13318_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16474__B1 _16219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18969_ _18969_/A VGND VGND VPWR VPWR _18982_/A sky130_fd_sc_hd__inv_2
XFILLER_100_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19412__B1 _19366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21980_ _21980_/A _21979_/X VGND VGND VPWR VPWR _21980_/X sky130_fd_sc_hd__or2_4
X_20931_ _20931_/A VGND VGND VPWR VPWR _20931_/X sky130_fd_sc_hd__buf_2
XFILLER_66_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16777__A1 _24404_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20862_ _16294_/Y _21093_/B _20856_/A _20861_/X VGND VGND VPWR VPWR _20863_/C sky130_fd_sc_hd__a211o_4
XFILLER_54_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23650_ _24823_/CLK _23650_/D HRESETn VGND VGND VPWR VPWR _23650_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23945__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19715__B2 _19710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22601_ _21434_/A VGND VGND VPWR VPWR _22601_/X sky130_fd_sc_hd__buf_2
X_20793_ _22953_/B _20792_/X VGND VGND VPWR VPWR _20794_/C sky130_fd_sc_hd__or2_4
XFILLER_81_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25169__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23581_ _23457_/CLK _23581_/D VGND VGND VPWR VPWR _17750_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13351__A _13338_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22532_ _20495_/A _22530_/X _20635_/C _22531_/X VGND VGND VPWR VPWR _22532_/X sky130_fd_sc_hd__a2bb2o_4
X_22463_ _22463_/A _20787_/B VGND VGND VPWR VPWR _22463_/X sky130_fd_sc_hd__or2_4
X_24202_ _24201_/CLK _16444_/X HRESETn VGND VGND VPWR VPWR _16443_/A sky130_fd_sc_hd__dfrtp_4
X_21414_ _24432_/Q _21710_/B VGND VGND VPWR VPWR _21414_/X sky130_fd_sc_hd__or2_4
X_22394_ _22306_/A _22384_/X _22387_/X _22394_/D VGND VGND VPWR VPWR _22394_/X sky130_fd_sc_hd__or4_4
X_25182_ _24847_/CLK _25182_/D HRESETn VGND VGND VPWR VPWR _11769_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18151__B1 _16063_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21345_ _21159_/A _19658_/Y VGND VGND VPWR VPWR _21345_/X sky130_fd_sc_hd__or2_4
XANTENNA__23027__A1 _21864_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24133_ _24101_/CLK _24133_/D HRESETn VGND VGND VPWR VPWR _24133_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16701__B2 _16700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21276_ _21276_/A VGND VGND VPWR VPWR _22351_/A sky130_fd_sc_hd__buf_2
XFILLER_116_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24064_ _24064_/CLK _24064_/D HRESETn VGND VGND VPWR VPWR _24064_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21589__A1 _12001_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11526__B1 _11525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20912__A _22014_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24733__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_HCLK clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_20227_ _20227_/A _20226_/X VGND VGND VPWR VPWR _20227_/X sky130_fd_sc_hd__or2_4
XANTENNA__22830__C _22830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17493__A _22395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23015_ _22982_/A _23012_/X _23013_/X _23015_/D VGND VGND VPWR VPWR _23015_/X sky130_fd_sc_hd__or4_4
XFILLER_131_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16723__A2_N _17614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23645__D sda_i_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20158_ _20158_/A VGND VGND VPWR VPWR _20158_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19403__B1 _19311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12980_ _12815_/Y _12984_/A _12805_/Y _12992_/B VGND VGND VPWR VPWR _12980_/X sky130_fd_sc_hd__or4_4
X_20089_ _20076_/Y VGND VGND VPWR VPWR _20089_/X sky130_fd_sc_hd__buf_2
X_24966_ _24587_/CLK _13520_/X HRESETn VGND VGND VPWR VPWR _20740_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_134_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16217__B1 _16216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11931_ _11919_/A VGND VGND VPWR VPWR _11931_/X sky130_fd_sc_hd__buf_2
X_23917_ _23908_/CLK _17994_/X HRESETn VGND VGND VPWR VPWR _23917_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16768__A1 _24403_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24897_ _24897_/CLK _13919_/X HRESETn VGND VGND VPWR VPWR _13830_/C sky130_fd_sc_hd__dfrtp_4
XANTENNA__16738__A2_N _17502_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15741__A _11944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14650_ _24726_/Q _14627_/X _24726_/Q _14627_/X VGND VGND VPWR VPWR _14651_/A sky130_fd_sc_hd__a2bb2o_4
X_11862_ _13053_/A VGND VGND VPWR VPWR _11862_/Y sky130_fd_sc_hd__inv_2
X_23848_ _23845_/CLK _23848_/D HRESETn VGND VGND VPWR VPWR _18211_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_45_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16280__A1_N _14897_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23686__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13601_ _13557_/B _13600_/Y _13594_/X _13586_/X _11663_/A VGND VGND VPWR VPWR _24950_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19706__B2 _19688_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14581_ _14581_/A VGND VGND VPWR VPWR _14581_/Y sky130_fd_sc_hd__inv_2
X_11793_ _11793_/A VGND VGND VPWR VPWR _11793_/Y sky130_fd_sc_hd__inv_2
X_23779_ _23668_/CLK _23779_/D HRESETn VGND VGND VPWR VPWR _23779_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22710__B1 _24416_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23615__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16320_ _16320_/A VGND VGND VPWR VPWR _16320_/Y sky130_fd_sc_hd__inv_2
X_13532_ _13532_/A _13532_/B VGND VGND VPWR VPWR _13533_/B sky130_fd_sc_hd__or2_4
XANTENNA__18390__B1 _24211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22574__A _14722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16251_ HWDATA[24] VGND VGND VPWR VPWR _16251_/X sky130_fd_sc_hd__buf_2
X_13463_ _13463_/A VGND VGND VPWR VPWR _13463_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16295__A1_N _16294_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15202_ _15208_/A _15211_/B VGND VGND VPWR VPWR _15203_/B sky130_fd_sc_hd__or2_4
X_12414_ _12409_/X _12414_/B VGND VGND VPWR VPWR _12415_/D sky130_fd_sc_hd__or2_4
XANTENNA__21277__B1 _22351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16182_ _16181_/Y _16178_/X _16087_/X _16178_/X VGND VGND VPWR VPWR _24304_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14951__B1 _14950_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13394_ _13381_/Y _13393_/Y SCLK_S2 _13392_/X VGND VGND VPWR VPWR _13394_/X sky130_fd_sc_hd__o22a_4
XFILLER_126_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_153_0_HCLK clkbuf_7_76_0_HCLK/X VGND VGND VPWR VPWR _25034_/CLK sky130_fd_sc_hd__clkbuf_1
X_15133_ _15154_/A _15131_/X _15133_/C VGND VGND VPWR VPWR _24679_/D sky130_fd_sc_hd__and3_4
XANTENNA__23018__A1 _24156_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12345_ _12344_/Y VGND VGND VPWR VPWR _12345_/X sky130_fd_sc_hd__buf_2
XFILLER_126_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15064_ _15064_/A _15064_/B VGND VGND VPWR VPWR _15065_/C sky130_fd_sc_hd__or2_4
X_19941_ _19941_/A VGND VGND VPWR VPWR _19941_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21918__A _20980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12276_ _12261_/A _12276_/B _12275_/Y VGND VGND VPWR VPWR _25112_/D sky130_fd_sc_hd__and3_4
XFILLER_107_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24474__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14015_ _14015_/A VGND VGND VPWR VPWR _14016_/A sky130_fd_sc_hd__buf_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15916__A _15916_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19872_ _21683_/B _19869_/X _19825_/X _19869_/X VGND VGND VPWR VPWR _23179_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24403__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16456__B1 _16455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18823_ _16291_/A VGND VGND VPWR VPWR _18823_/X sky130_fd_sc_hd__buf_2
XFILLER_7_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22529__B1 _13335_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15966_ _15987_/A VGND VGND VPWR VPWR _15966_/X sky130_fd_sc_hd__buf_2
X_18754_ _18754_/A VGND VGND VPWR VPWR _18754_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17405__C1 _17336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14917_ _14915_/A _24262_/Q _15108_/C _14916_/Y VGND VGND VPWR VPWR _14918_/D sky130_fd_sc_hd__o22a_4
X_17705_ _15712_/X _15713_/X _13474_/A _15813_/X VGND VGND VPWR VPWR _17705_/X sky130_fd_sc_hd__a211o_4
X_15897_ _16376_/A VGND VGND VPWR VPWR _15897_/X sky130_fd_sc_hd__buf_2
X_18685_ _16216_/A VGND VGND VPWR VPWR _18685_/X sky130_fd_sc_hd__buf_2
X_14848_ _14842_/X _14843_/X _14845_/X _14847_/X VGND VGND VPWR VPWR _14848_/X sky130_fd_sc_hd__or4_4
X_17636_ _17636_/A VGND VGND VPWR VPWR _17636_/X sky130_fd_sc_hd__buf_2
X_17567_ _17547_/X _17563_/B _17566_/X VGND VGND VPWR VPWR _17567_/X sky130_fd_sc_hd__and3_4
X_14779_ _24113_/Q VGND VGND VPWR VPWR _14779_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14267__A _13619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22701__B1 _12088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16518_ _16499_/A VGND VGND VPWR VPWR _16518_/X sky130_fd_sc_hd__buf_2
X_19306_ _19302_/Y _19305_/X _19170_/X _19305_/X VGND VGND VPWR VPWR _23382_/D sky130_fd_sc_hd__a2bb2o_4
X_17498_ _17498_/A VGND VGND VPWR VPWR _17498_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16449_ _16448_/Y _16446_/X _16279_/X _16446_/X VGND VGND VPWR VPWR _24200_/D sky130_fd_sc_hd__a2bb2o_4
X_19237_ _18018_/X _19282_/B _19236_/X VGND VGND VPWR VPWR _19238_/A sky130_fd_sc_hd__or3_4
XFILLER_121_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19168_ _19167_/X VGND VGND VPWR VPWR _19175_/A sky130_fd_sc_hd__inv_2
XANTENNA__14942__B1 _14941_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18119_ _18117_/Y _18113_/X _18120_/A _18118_/X VGND VGND VPWR VPWR _18119_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23009__A1 _16621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15098__A _15158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19099_ _23454_/Q VGND VGND VPWR VPWR _19099_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23009__B2 _21694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21130_ _21130_/A VGND VGND VPWR VPWR _21130_/X sky130_fd_sc_hd__buf_2
XFILLER_132_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21828__A _20980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21061_ _21040_/X _21049_/Y _22245_/A _21060_/X VGND VGND VPWR VPWR _21061_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22001__A1_N _12408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24144__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20012_ _20012_/A VGND VGND VPWR VPWR _22092_/B sky130_fd_sc_hd__inv_2
XANTENNA__16447__B1 _16100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24820_ _24823_/CLK _14210_/X HRESETn VGND VGND VPWR VPWR _20193_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_39_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12484__A1 _12474_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24751_ _25009_/CLK _24751_/D HRESETn VGND VGND VPWR VPWR _14430_/A sky130_fd_sc_hd__dfrtp_4
X_21963_ _21214_/A _19513_/Y _21202_/A VGND VGND VPWR VPWR _21963_/X sky130_fd_sc_hd__o21a_4
X_23702_ _23702_/CLK _23702_/D HRESETn VGND VGND VPWR VPWR _13506_/A sky130_fd_sc_hd__dfrtp_4
X_20914_ _21591_/B VGND VGND VPWR VPWR _22154_/B sky130_fd_sc_hd__buf_2
XFILLER_82_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24682_ _24676_/CLK _15097_/X HRESETn VGND VGND VPWR VPWR _15096_/A sky130_fd_sc_hd__dfrtp_4
X_21894_ _14270_/Y _21544_/A _24790_/Q _21180_/X VGND VGND VPWR VPWR _21894_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16094__A2_N _16090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23633_ _23641_/CLK _23633_/D HRESETn VGND VGND VPWR VPWR _20292_/A sky130_fd_sc_hd__dfrtp_4
X_20845_ _20719_/A _14015_/A _23657_/Q _21088_/A VGND VGND VPWR VPWR _20849_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13081__A _11751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23564_ _23563_/CLK _18791_/X VGND VGND VPWR VPWR _23564_/Q sky130_fd_sc_hd__dfxtp_4
X_20776_ _22438_/A VGND VGND VPWR VPWR _22971_/A sky130_fd_sc_hd__buf_2
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20907__A _20833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22515_ _24483_/Q _22757_/B VGND VGND VPWR VPWR _22515_/X sky130_fd_sc_hd__or2_4
XANTENNA__17488__A _20778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23495_ _23128_/CLK _18987_/X VGND VGND VPWR VPWR _18986_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24985__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20626__B _13537_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22446_ _24269_/Q _22227_/B _22435_/X _22445_/X VGND VGND VPWR VPWR _22446_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24914__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25165_ _23898_/CLK _25165_/D HRESETn VGND VGND VPWR VPWR _11871_/B sky130_fd_sc_hd__dfrtp_4
X_22377_ _22377_/A _22527_/B VGND VGND VPWR VPWR _22377_/X sky130_fd_sc_hd__and2_4
XFILLER_100_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19872__B1 _19825_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_226_0_HCLK clkbuf_8_227_0_HCLK/A VGND VGND VPWR VPWR _24307_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_108_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12130_ _12237_/A _24559_/Q _12237_/A _24559_/Q VGND VGND VPWR VPWR _12130_/X sky130_fd_sc_hd__a2bb2o_4
X_24116_ _24112_/CLK _16637_/X HRESETn VGND VGND VPWR VPWR _24116_/Q sky130_fd_sc_hd__dfrtp_4
X_21328_ _21169_/A _21328_/B VGND VGND VPWR VPWR _21328_/X sky130_fd_sc_hd__or2_4
XFILLER_123_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25096_ _25097_/CLK _25096_/D HRESETn VGND VGND VPWR VPWR _12317_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12361__A2_N _22373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12061_ _13612_/A _12061_/B _24618_/Q VGND VGND VPWR VPWR _12062_/A sky130_fd_sc_hd__or3_4
X_21259_ _21259_/A VGND VGND VPWR VPWR _21259_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15736__A _15741_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24047_ _24604_/CLK _17103_/Y HRESETn VGND VGND VPWR VPWR _24047_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21457__B _21457_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18112__A _18112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21982__A1 _21178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15820_ _22933_/B VGND VGND VPWR VPWR _15824_/A sky130_fd_sc_hd__buf_2
XANTENNA__21982__B2 _16393_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23867__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15751_ _15750_/Y VGND VGND VPWR VPWR _15757_/A sky130_fd_sc_hd__buf_2
XANTENNA__21473__A _21339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12963_ _12963_/A _12933_/D VGND VGND VPWR VPWR _12964_/B sky130_fd_sc_hd__or2_4
XFILLER_57_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12475__A1 _12412_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24949_ _23925_/CLK _13603_/X HRESETn VGND VGND VPWR VPWR _11687_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_92_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13672__B1 _13635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21734__B2 _21179_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14702_ _24707_/Q VGND VGND VPWR VPWR _14702_/Y sky130_fd_sc_hd__inv_2
X_11914_ _23789_/Q _11905_/X _11911_/Y VGND VGND VPWR VPWR _11914_/X sky130_fd_sc_hd__o21a_4
X_18470_ _18470_/A _18470_/B VGND VGND VPWR VPWR _18470_/X sky130_fd_sc_hd__or2_4
XANTENNA__18485__C _18485_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15682_ _12326_/Y _15680_/X _11570_/X _15680_/X VGND VGND VPWR VPWR _24485_/D sky130_fd_sc_hd__a2bb2o_4
X_12894_ _12894_/A _12894_/B VGND VGND VPWR VPWR _12894_/X sky130_fd_sc_hd__or2_4
XFILLER_61_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17421_ _17423_/A _17421_/B _17420_/Y VGND VGND VPWR VPWR _23987_/D sky130_fd_sc_hd__and3_4
X_14633_ _14633_/A VGND VGND VPWR VPWR _14633_/X sky130_fd_sc_hd__buf_2
XFILLER_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11845_ _11843_/Y _11840_/X _11844_/X _11840_/X VGND VGND VPWR VPWR _25173_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17352_ _17352_/A _17352_/B VGND VGND VPWR VPWR _17354_/B sky130_fd_sc_hd__or2_4
XFILLER_57_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14564_ _17947_/A VGND VGND VPWR VPWR _14564_/X sky130_fd_sc_hd__buf_2
X_11776_ _25178_/Q _11776_/B VGND VGND VPWR VPWR _11817_/A sky130_fd_sc_hd__and2_4
X_16303_ _18258_/A _16302_/Y _16219_/X _16302_/Y VGND VGND VPWR VPWR _16303_/X sky130_fd_sc_hd__a2bb2o_4
X_13515_ _20542_/A _20542_/B _20545_/A _13514_/X VGND VGND VPWR VPWR _13515_/X sky130_fd_sc_hd__or4_4
XFILLER_53_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17283_ _11557_/Y _24000_/Q _25200_/Q _17415_/A VGND VGND VPWR VPWR _17283_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14495_ _14471_/A _14489_/X _14494_/X _14490_/Y VGND VGND VPWR VPWR _14495_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_6_36_0_HCLK clkbuf_6_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_73_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19022_ _23482_/Q VGND VGND VPWR VPWR _21505_/B sky130_fd_sc_hd__inv_2
X_16234_ _16234_/A VGND VGND VPWR VPWR _16234_/X sky130_fd_sc_hd__buf_2
XFILLER_70_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13446_ _13446_/A VGND VGND VPWR VPWR _13446_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24655__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18006__B _11944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16165_ _16165_/A VGND VGND VPWR VPWR _16165_/X sky130_fd_sc_hd__buf_2
X_13377_ _13363_/A VGND VGND VPWR VPWR _13377_/X sky130_fd_sc_hd__buf_2
XANTENNA__12335__A _24474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15116_ _15138_/A _15138_/B _15103_/X _15115_/X VGND VGND VPWR VPWR _15117_/C sky130_fd_sc_hd__or4_4
X_12328_ _12328_/A VGND VGND VPWR VPWR _12328_/Y sky130_fd_sc_hd__inv_2
X_16096_ _16096_/A VGND VGND VPWR VPWR _16096_/X sky130_fd_sc_hd__buf_2
XFILLER_5_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15047_ _15042_/A _15019_/X _15027_/X _15044_/B VGND VGND VPWR VPWR _15047_/X sky130_fd_sc_hd__a211o_4
X_19924_ _23158_/Q VGND VGND VPWR VPWR _22064_/B sky130_fd_sc_hd__inv_2
X_12259_ _25115_/Q _12259_/B VGND VGND VPWR VPWR _12261_/B sky130_fd_sc_hd__or2_4
XFILLER_68_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16429__B1 _16264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19855_ _19853_/Y _19854_/X _19832_/X _19854_/X VGND VGND VPWR VPWR _19855_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18806_ _13038_/B VGND VGND VPWR VPWR _18806_/Y sky130_fd_sc_hd__inv_2
X_19786_ _19780_/Y VGND VGND VPWR VPWR _19786_/X sky130_fd_sc_hd__buf_2
X_16998_ _16183_/Y _24041_/Q _16183_/Y _24041_/Q VGND VGND VPWR VPWR _16998_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21383__A _21383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18737_ _18732_/Y _18736_/X _17199_/X _18736_/X VGND VGND VPWR VPWR _23582_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15949_ _15947_/Y _15948_/X _15855_/X _15948_/X VGND VGND VPWR VPWR _24381_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21725__B2 _21570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15381__A _15358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18668_ _18682_/A VGND VGND VPWR VPWR _18668_/X sky130_fd_sc_hd__buf_2
XFILLER_64_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17619_ _17619_/A _17615_/X _17618_/Y VGND VGND VPWR VPWR _23944_/D sky130_fd_sc_hd__and3_4
XFILLER_52_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_118_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_237_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18599_ _16304_/Y _18442_/A _16304_/Y _18442_/A VGND VGND VPWR VPWR _18599_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21489__B1 _20820_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20630_ _20635_/A VGND VGND VPWR VPWR _20630_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11523__A2_N _11521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18354__B1 _24217_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20727__A _23666_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20561_ _20560_/X VGND VGND VPWR VPWR _20561_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20700__A2 _23616_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22300_ _24300_/Q _22246_/B VGND VGND VPWR VPWR _22300_/X sky130_fd_sc_hd__or2_4
XFILLER_137_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20492_ _20495_/A _20495_/B _20491_/X VGND VGND VPWR VPWR _20492_/X sky130_fd_sc_hd__o21a_4
XFILLER_30_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23280_ _23303_/CLK _23280_/D VGND VGND VPWR VPWR _19590_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_121_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24396__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22989__B1 _22858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22231_ _22551_/A VGND VGND VPWR VPWR _22231_/X sky130_fd_sc_hd__buf_2
XANTENNA__22453__A2 _21576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24325__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16668__B1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22162_ _24510_/Q _21047_/X _20744_/X _22161_/X VGND VGND VPWR VPWR _22162_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16132__A2 _16135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21113_ _21097_/B _21113_/B _21113_/C _21275_/A VGND VGND VPWR VPWR _21113_/X sky130_fd_sc_hd__or4_4
X_22093_ _22089_/A _22091_/X _22092_/X VGND VGND VPWR VPWR _22093_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_56_0_HCLK clkbuf_7_28_0_HCLK/X VGND VGND VPWR VPWR _24008_/CLK sky130_fd_sc_hd__clkbuf_1
X_21044_ _21044_/A _21043_/X VGND VGND VPWR VPWR _21044_/X sky130_fd_sc_hd__or2_4
XFILLER_120_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23807__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21964__A1 _21224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12411__C _12410_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23960__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24803_ _24811_/CLK _14258_/X HRESETn VGND VGND VPWR VPWR _14257_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__25184__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13654__B1 _11594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22995_ _22429_/B _22991_/X _22407_/X _22994_/X VGND VGND VPWR VPWR _22995_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15291__A _14218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24734_ _23568_/CLK _24734_/D HRESETn VGND VGND VPWR VPWR _14581_/A sky130_fd_sc_hd__dfrtp_4
X_21946_ _21367_/A _21946_/B VGND VGND VPWR VPWR _21946_/X sky130_fd_sc_hd__or2_4
XFILLER_76_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25113__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24665_ _24671_/CLK _15183_/X HRESETn VGND VGND VPWR VPWR _24665_/Q sky130_fd_sc_hd__dfrtp_4
X_21877_ _19263_/A _21082_/B _15428_/X _21876_/X VGND VGND VPWR VPWR _21877_/X sky130_fd_sc_hd__a211o_4
XPHY_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11630_/A VGND VGND VPWR VPWR _15282_/A sky130_fd_sc_hd__buf_2
XPHY_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23616_ _23774_/CLK _23616_/D HRESETn VGND VGND VPWR VPWR _23616_/Q sky130_fd_sc_hd__dfrtp_4
X_20828_ _24462_/Q _20826_/X _20738_/B _20827_/X VGND VGND VPWR VPWR _20828_/X sky130_fd_sc_hd__o22a_4
XPHY_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22141__A1 _11992_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24596_ _24596_/CLK _15375_/X HRESETn VGND VGND VPWR VPWR _15373_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _11533_/X _11535_/X HWDATA[21] _25211_/Q _11537_/X VGND VGND VPWR VPWR _11561_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23547_ _23482_/CLK _18841_/X VGND VGND VPWR VPWR _23547_/Q sky130_fd_sc_hd__dfxtp_4
X_20759_ _20758_/X VGND VGND VPWR VPWR _20759_/X sky130_fd_sc_hd__buf_2
XANTENNA__18896__B2 _18876_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13300_ _13300_/A _13300_/B VGND VGND VPWR VPWR _13302_/B sky130_fd_sc_hd__or2_4
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14280_ _14273_/A VGND VGND VPWR VPWR _14280_/X sky130_fd_sc_hd__buf_2
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23478_ _23537_/CLK _19036_/X VGND VGND VPWR VPWR _13022_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ _13159_/X _13231_/B _13231_/C VGND VGND VPWR VPWR _13231_/X sky130_fd_sc_hd__and3_4
XFILLER_10_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25217_ _25217_/CLK _25217_/D HRESETn VGND VGND VPWR VPWR _25217_/Q sky130_fd_sc_hd__dfrtp_4
X_22429_ _24041_/Q _22429_/B VGND VGND VPWR VPWR _22433_/B sky130_fd_sc_hd__or2_4
XANTENNA__24066__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13162_ _13230_/A _23131_/Q VGND VGND VPWR VPWR _13162_/X sky130_fd_sc_hd__or2_4
XANTENNA__21652__B1 _21642_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21468__A _21144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25148_ _24824_/CLK _25148_/D HRESETn VGND VGND VPWR VPWR _11983_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_124_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12113_ _12113_/A VGND VGND VPWR VPWR _12265_/B sky130_fd_sc_hd__inv_2
X_13093_ _13169_/A VGND VGND VPWR VPWR _13137_/A sky130_fd_sc_hd__buf_2
X_17970_ _16022_/Y _17970_/B _17970_/C VGND VGND VPWR VPWR _17970_/X sky130_fd_sc_hd__and3_4
XANTENNA__16674__A3 _16558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25079_ _25090_/CLK _25079_/D HRESETn VGND VGND VPWR VPWR _12344_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_3_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21404__B1 _21256_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12044_ _11985_/Y _12043_/X _11985_/Y _12043_/X VGND VGND VPWR VPWR _12044_/X sky130_fd_sc_hd__a2bb2o_4
X_16921_ _16832_/Y _16778_/Y _16921_/C _16921_/D VGND VGND VPWR VPWR _16922_/B sky130_fd_sc_hd__or4_4
XFILLER_133_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19640_ _19640_/A VGND VGND VPWR VPWR _20964_/B sky130_fd_sc_hd__inv_2
XFILLER_120_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16852_ _16879_/A _16852_/B VGND VGND VPWR VPWR _16853_/B sky130_fd_sc_hd__or2_4
XFILLER_78_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15803_ _12826_/Y _15757_/A _15709_/X _15757_/A VGND VGND VPWR VPWR _15803_/X sky130_fd_sc_hd__a2bb2o_4
X_16783_ _16756_/X _16764_/X _16783_/C _16783_/D VGND VGND VPWR VPWR _16811_/A sky130_fd_sc_hd__or4_4
X_19571_ _23287_/Q VGND VGND VPWR VPWR _19571_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15913__B _15418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13995_ _13938_/X _13994_/Y _24811_/Q _13938_/X VGND VGND VPWR VPWR _24883_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23630__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15734_ _15716_/A _15733_/X _15726_/A VGND VGND VPWR VPWR _24464_/D sky130_fd_sc_hd__o21a_4
X_18522_ _18448_/A VGND VGND VPWR VPWR _18540_/A sky130_fd_sc_hd__buf_2
X_12946_ _12943_/C _12943_/D VGND VGND VPWR VPWR _12947_/B sky130_fd_sc_hd__or2_4
XFILLER_4_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18584__B1 _24243_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15665_ _15695_/A VGND VGND VPWR VPWR _15666_/A sky130_fd_sc_hd__buf_2
X_18453_ _18453_/A VGND VGND VPWR VPWR _18453_/Y sky130_fd_sc_hd__inv_2
X_12877_ _12815_/Y _12984_/A _12863_/Y _12876_/X VGND VGND VPWR VPWR _12974_/A sky130_fd_sc_hd__or4_4
X_14616_ _24730_/Q VGND VGND VPWR VPWR _14617_/C sky130_fd_sc_hd__inv_2
X_17404_ _17423_/A _17402_/X _17404_/C VGND VGND VPWR VPWR _17404_/X sky130_fd_sc_hd__and3_4
X_11828_ _11780_/Y _11828_/B _11694_/X VGND VGND VPWR VPWR _11828_/X sky130_fd_sc_hd__or3_4
X_18384_ _16443_/Y _23825_/Q _16443_/Y _23825_/Q VGND VGND VPWR VPWR _18384_/X sky130_fd_sc_hd__a2bb2o_4
X_15596_ HWDATA[25] VGND VGND VPWR VPWR _15596_/X sky130_fd_sc_hd__buf_2
XANTENNA__24836__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17300_/X VGND VGND VPWR VPWR _17622_/B sky130_fd_sc_hd__inv_2
XPHY_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14482_/X _14491_/X _19883_/B _14437_/X VGND VGND VPWR VPWR _14547_/X sky130_fd_sc_hd__o22a_4
X_11759_ _13050_/A _11758_/X _13050_/A _11758_/X VGND VGND VPWR VPWR _11759_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22683__A2 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17266_ _23996_/Q VGND VGND VPWR VPWR _17266_/Y sky130_fd_sc_hd__inv_2
X_14478_ _14476_/Y _14482_/A VGND VGND VPWR VPWR _14479_/A sky130_fd_sc_hd__or2_4
XFILLER_31_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16217_ _16215_/Y _16138_/A _16216_/X _16138_/A VGND VGND VPWR VPWR _16217_/X sky130_fd_sc_hd__a2bb2o_4
X_19005_ _19005_/A VGND VGND VPWR VPWR _19005_/Y sky130_fd_sc_hd__inv_2
X_13429_ _14414_/A VGND VGND VPWR VPWR _13429_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17197_ _13619_/X _17197_/B VGND VGND VPWR VPWR _17213_/A sky130_fd_sc_hd__nor2_4
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19836__B1 _19835_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16148_ _16147_/Y _16145_/X _15837_/X _16145_/X VGND VGND VPWR VPWR _24317_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_6_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16079_ _16078_/Y _16076_/X _15775_/X _16076_/X VGND VGND VPWR VPWR _24342_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21097__B _21097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22199__A1 _22195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22199__B2 _22198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23789__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19907_ _22079_/B _19906_/X _19815_/X _19906_/X VGND VGND VPWR VPWR _19907_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23718__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17591__A _22307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19838_ _19837_/Y _19831_/X _19506_/X _19831_/A VGND VGND VPWR VPWR _23191_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23780__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19769_ _19769_/A VGND VGND VPWR VPWR _21463_/B sky130_fd_sc_hd__inv_2
XFILLER_83_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13636__B1 _13635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22002__A _21245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21800_ _21799_/A _20070_/A VGND VGND VPWR VPWR _21800_/X sky130_fd_sc_hd__or2_4
X_22780_ _24526_/Q _20799_/X _20801_/X _22779_/X VGND VGND VPWR VPWR _22781_/C sky130_fd_sc_hd__a211o_4
XANTENNA__22371__A1 _22369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21731_ _20819_/X _21727_/X _22407_/A _21730_/X VGND VGND VPWR VPWR _21731_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21841__A _15456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19311__A _18743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24450_ _24459_/CLK _15769_/X HRESETn VGND VGND VPWR VPWR _22703_/A sky130_fd_sc_hd__dfrtp_4
X_21662_ _14529_/X VGND VGND VPWR VPWR _21665_/A sky130_fd_sc_hd__buf_2
XFILLER_52_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14061__B1 _13638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24577__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23401_ _23401_/CLK _19252_/X VGND VGND VPWR VPWR _19250_/A sky130_fd_sc_hd__dfxtp_4
X_20613_ _20598_/X _20612_/X _24170_/Q _20603_/X VGND VGND VPWR VPWR _20613_/X sky130_fd_sc_hd__a2bb2o_4
X_24381_ _24378_/CLK _24381_/D HRESETn VGND VGND VPWR VPWR _22706_/A sky130_fd_sc_hd__dfrtp_4
X_21593_ _16464_/Y _22840_/A _16300_/A _21592_/X VGND VGND VPWR VPWR _21600_/C sky130_fd_sc_hd__a211o_4
XANTENNA__24506__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23332_ _23332_/CLK _23332_/D VGND VGND VPWR VPWR _19447_/A sky130_fd_sc_hd__dfxtp_4
X_20544_ _20419_/X _20543_/X _15329_/A _20465_/X VGND VGND VPWR VPWR _20544_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22426__A2 _20799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23263_ _23356_/CLK _19642_/X VGND VGND VPWR VPWR _19640_/A sky130_fd_sc_hd__dfxtp_4
X_20475_ _20472_/Y _20473_/Y _20474_/X VGND VGND VPWR VPWR _20475_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22391__B _22999_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12375__B1 _12489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25002_ _25002_/CLK _25002_/D HRESETn VGND VGND VPWR VPWR _25002_/Q sky130_fd_sc_hd__dfrtp_4
X_22214_ _22214_/A _21357_/X VGND VGND VPWR VPWR _22214_/X sky130_fd_sc_hd__and2_4
XFILLER_10_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23194_ _23154_/CLK _19829_/X VGND VGND VPWR VPWR _23194_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_134_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15286__A _15801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22145_ _21570_/X VGND VGND VPWR VPWR _22879_/A sky130_fd_sc_hd__buf_2
XANTENNA__15313__B1 HADDR[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22076_ _21786_/A _19573_/Y VGND VGND VPWR VPWR _22076_/X sky130_fd_sc_hd__or2_4
XFILLER_82_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13518__B _13517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21027_ _21027_/A VGND VGND VPWR VPWR _21027_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12800_ _22161_/A VGND VGND VPWR VPWR _12800_/Y sky130_fd_sc_hd__inv_2
X_13780_ _13770_/A _13780_/B _13773_/D VGND VGND VPWR VPWR _13795_/A sky130_fd_sc_hd__or3_4
X_22978_ _22919_/A _22978_/B _22971_/X _22977_/X VGND VGND VPWR VPWR _22978_/X sky130_fd_sc_hd__or4_4
XANTENNA__22362__A1 _22116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22362__B2 _22118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12731_ _12731_/A _12728_/X VGND VGND VPWR VPWR _12732_/C sky130_fd_sc_hd__or2_4
X_24717_ _23664_/CLK _24717_/D HRESETn VGND VGND VPWR VPWR _14609_/A sky130_fd_sc_hd__dfrtp_4
X_21929_ _21155_/A _21927_/X _21928_/X VGND VGND VPWR VPWR _21929_/X sky130_fd_sc_hd__and3_4
XFILLER_43_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16845__A _16846_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15450_ _14432_/X _15441_/B VGND VGND VPWR VPWR _15450_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__19221__A _11625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12662_ _12727_/A _12915_/C VGND VGND VPWR VPWR _12663_/B sky130_fd_sc_hd__and2_4
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24648_ _24643_/CLK _24648_/D HRESETn VGND VGND VPWR VPWR _13753_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_71_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_101_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_203_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14386_/A _14399_/X _14400_/Y _13608_/X _13416_/A VGND VGND VPWR VPWR _24764_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11609_/Y _11610_/X _11612_/X _11610_/X VGND VGND VPWR VPWR _11613_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11989__A _15271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15358_/X VGND VGND VPWR VPWR _15381_/X sky130_fd_sc_hd__buf_2
XFILLER_106_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _12593_/A VGND VGND VPWR VPWR _12593_/Y sky130_fd_sc_hd__inv_2
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24579_ _25183_/CLK _24579_/D HRESETn VGND VGND VPWR VPWR _14433_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14365__A HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24247__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17120_ _17101_/A _17118_/X _17120_/C VGND VGND VPWR VPWR _24042_/D sky130_fd_sc_hd__and3_4
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ _14329_/A _14330_/X _14286_/A _14331_/X VGND VGND VPWR VPWR _24779_/D sky130_fd_sc_hd__o22a_4
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11544_ _25216_/Q VGND VGND VPWR VPWR _11544_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_5_21_0_HCLK_A clkbuf_4_10_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17051_ _24058_/Q _17051_/B VGND VGND VPWR VPWR _17051_/Y sky130_fd_sc_hd__nand2_4
XFILLER_7_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ _14262_/Y _14260_/X _14094_/X _14260_/X VGND VGND VPWR VPWR _24801_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17676__A _17918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16002_ _16001_/Y _15922_/X _15291_/X _15922_/X VGND VGND VPWR VPWR _16002_/X sky130_fd_sc_hd__a2bb2o_4
X_13214_ _13278_/A _13212_/X _13213_/X VGND VGND VPWR VPWR _13214_/X sky130_fd_sc_hd__and3_4
XFILLER_13_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14194_ _11512_/Y VGND VGND VPWR VPWR _14195_/C sky130_fd_sc_hd__buf_2
XFILLER_125_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19294__B2 _19289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13145_ _13169_/A VGND VGND VPWR VPWR _13146_/A sky130_fd_sc_hd__buf_2
XFILLER_124_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23882__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13076_ _13076_/A VGND VGND VPWR VPWR _13127_/A sky130_fd_sc_hd__buf_2
X_17953_ _17889_/A _17951_/X _17952_/X VGND VGND VPWR VPWR _17954_/C sky130_fd_sc_hd__and3_4
XFILLER_2_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12027_ _12026_/X VGND VGND VPWR VPWR _12027_/Y sky130_fd_sc_hd__inv_2
X_16904_ _16823_/Y _16898_/B VGND VGND VPWR VPWR _16904_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22050__B1 _20820_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25035__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17884_ _17816_/A _17884_/B VGND VGND VPWR VPWR _17886_/B sky130_fd_sc_hd__or2_4
X_19623_ _19623_/A VGND VGND VPWR VPWR _19636_/A sky130_fd_sc_hd__inv_2
XFILLER_38_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16835_ _16835_/A VGND VGND VPWR VPWR _16922_/A sky130_fd_sc_hd__inv_2
XFILLER_47_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19554_ _19554_/A VGND VGND VPWR VPWR _19554_/Y sky130_fd_sc_hd__inv_2
X_13978_ _13956_/X _13977_/X _24800_/Q _13963_/X VGND VGND VPWR VPWR _13978_/Y sky130_fd_sc_hd__a22oi_4
X_16766_ _24414_/Q _16765_/A _15859_/Y _16765_/Y VGND VGND VPWR VPWR _16766_/X sky130_fd_sc_hd__o22a_4
XFILLER_93_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14291__B1 _14232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18505_ _18434_/D _18495_/D _18475_/X _18503_/B VGND VGND VPWR VPWR _18506_/A sky130_fd_sc_hd__a211o_4
X_12929_ _12952_/A _12917_/B _12929_/C VGND VGND VPWR VPWR _12929_/X sky130_fd_sc_hd__and3_4
X_15717_ _15717_/A _15717_/B _15717_/C VGND VGND VPWR VPWR _15717_/X sky130_fd_sc_hd__or3_4
X_16697_ _23960_/Q VGND VGND VPWR VPWR _16697_/Y sky130_fd_sc_hd__inv_2
X_19485_ _19484_/Y _19480_/X _19392_/X _19467_/Y VGND VGND VPWR VPWR _23319_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22476__B _22473_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18436_ _18485_/D _18436_/B VGND VGND VPWR VPWR _18468_/B sky130_fd_sc_hd__or2_4
X_15648_ _15418_/A _15459_/A VGND VGND VPWR VPWR _15648_/X sky130_fd_sc_hd__or2_4
XFILLER_107_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24670__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15579_ _15578_/X VGND VGND VPWR VPWR _15741_/B sky130_fd_sc_hd__buf_2
X_18367_ _18359_/X _18362_/X _18364_/X _18366_/X VGND VGND VPWR VPWR _18367_/X sky130_fd_sc_hd__or4_4
XANTENNA__18970__A _18982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17318_ _17318_/A VGND VGND VPWR VPWR _17320_/A sky130_fd_sc_hd__inv_2
XFILLER_33_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18298_ _18298_/A VGND VGND VPWR VPWR _23857_/D sky130_fd_sc_hd__inv_2
XFILLER_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17249_ _11640_/Y _23978_/Q _11640_/Y _23978_/Q VGND VGND VPWR VPWR _17249_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16490__A _24184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20260_ _23767_/Q _20265_/B _20232_/X VGND VGND VPWR VPWR _20260_/X sky130_fd_sc_hd__a21o_4
XFILLER_115_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19285__B2 _19284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12130__A2_N _24559_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13619__A _16305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20191_ _13908_/A _20191_/B VGND VGND VPWR VPWR _20194_/C sky130_fd_sc_hd__and2_4
XFILLER_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23950_ _24079_/CLK _17603_/X HRESETn VGND VGND VPWR VPWR _16699_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21555__B _22227_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22592__A1 _22116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18796__B1 _18795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12145__A2_N _24549_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22592__B2 _22118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22901_ _12417_/A _22178_/A _24054_/Q _22652_/X VGND VGND VPWR VPWR _22904_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12775__A2_N _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23881_ _23885_/CLK _23881_/D HRESETn VGND VGND VPWR VPWR _23881_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_38_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17992__A1_N _11680_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22832_ _22832_/A _22813_/X _22832_/C _22831_/X VGND VGND VPWR VPWR HRDATA[25] sky130_fd_sc_hd__or4_4
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24758__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22763_ _22763_/A _22638_/X VGND VGND VPWR VPWR _22763_/X sky130_fd_sc_hd__or2_4
XFILLER_52_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24502_ _24502_/CLK _24502_/D HRESETn VGND VGND VPWR VPWR _20822_/A sky130_fd_sc_hd__dfrtp_4
X_21714_ _21713_/X VGND VGND VPWR VPWR _21857_/A sky130_fd_sc_hd__inv_2
XANTENNA__19041__A _18743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22694_ _24243_/Q _21553_/X _22148_/X _22693_/X VGND VGND VPWR VPWR _22694_/X sky130_fd_sc_hd__a211o_4
XFILLER_25_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24433_ _24372_/CLK _24433_/D HRESETn VGND VGND VPWR VPWR _15797_/A sky130_fd_sc_hd__dfrtp_4
X_21645_ _21648_/A _23105_/Q _18089_/A _20066_/Y VGND VGND VPWR VPWR _21645_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15782__B1 _22463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24340__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24364_ _24405_/CLK _15994_/X HRESETn VGND VGND VPWR VPWR _15991_/A sky130_fd_sc_hd__dfrtp_4
X_21576_ _21280_/A VGND VGND VPWR VPWR _21576_/X sky130_fd_sc_hd__buf_2
XANTENNA__18720__B1 _17205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23315_ _23313_/CLK _19497_/X VGND VGND VPWR VPWR _23315_/Q sky130_fd_sc_hd__dfxtp_4
X_20527_ _23720_/Q VGND VGND VPWR VPWR _20527_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17496__A _22434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24295_ _24319_/CLK _24295_/D HRESETn VGND VGND VPWR VPWR _16202_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_118_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23246_ _23246_/CLK _23246_/D VGND VGND VPWR VPWR _23246_/Q sky130_fd_sc_hd__dfxtp_4
X_20458_ _20457_/Y _20453_/Y _13506_/X VGND VGND VPWR VPWR _20458_/X sky130_fd_sc_hd__o21a_4
XFILLER_49_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23177_ _25112_/CLK _19877_/X VGND VGND VPWR VPWR _19875_/A sky130_fd_sc_hd__dfxtp_4
X_20389_ _20389_/A _20389_/B VGND VGND VPWR VPWR _20390_/B sky130_fd_sc_hd__nand2_4
XFILLER_97_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20830__A1 _21716_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22128_ _22127_/X VGND VGND VPWR VPWR _22128_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20830__B2 _22859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_26_0_HCLK clkbuf_7_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_53_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_14950_ _24665_/Q VGND VGND VPWR VPWR _14950_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15744__A _16305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22059_ _14487_/X _22059_/B _22058_/X VGND VGND VPWR VPWR _22059_/X sky130_fd_sc_hd__or3_4
XFILLER_0_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_89_0_HCLK clkbuf_6_44_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_89_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16559__B _16235_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13901_ _20251_/A _13896_/X _13900_/X _13866_/B _13893_/X VGND VGND VPWR VPWR _24909_/D
+ sky130_fd_sc_hd__a32o_4
X_14881_ _14881_/A _14995_/A VGND VGND VPWR VPWR _14881_/X sky130_fd_sc_hd__or2_4
XFILLER_29_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13832_ _13869_/D VGND VGND VPWR VPWR _13833_/D sky130_fd_sc_hd__inv_2
X_16620_ _15463_/A VGND VGND VPWR VPWR _16621_/A sky130_fd_sc_hd__buf_2
XANTENNA__24499__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16551_ _24160_/Q VGND VGND VPWR VPWR _16551_/Y sky130_fd_sc_hd__inv_2
X_13763_ _13763_/A VGND VGND VPWR VPWR _14071_/D sky130_fd_sc_hd__inv_2
XFILLER_95_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24428__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17211__B1 _16211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12714_ _12607_/Y _12714_/B VGND VGND VPWR VPWR _12714_/X sky130_fd_sc_hd__or2_4
X_15502_ _15482_/X _15483_/X _15501_/X _24558_/Q _15495_/X VGND VGND VPWR VPWR _24558_/D
+ sky130_fd_sc_hd__a32o_4
X_16482_ _16477_/Y _16481_/X _16141_/X _16481_/X VGND VGND VPWR VPWR _24188_/D sky130_fd_sc_hd__a2bb2o_4
X_19270_ _23394_/Q VGND VGND VPWR VPWR _21756_/B sky130_fd_sc_hd__buf_2
XFILLER_43_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13694_ _13678_/X _13692_/X _14077_/A _13693_/X VGND VGND VPWR VPWR _13694_/X sky130_fd_sc_hd__o22a_4
XFILLER_16_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15433_ _16302_/A _16475_/B VGND VGND VPWR VPWR _15433_/X sky130_fd_sc_hd__or2_4
X_18221_ _18221_/A _18198_/Y _18221_/C VGND VGND VPWR VPWR _18222_/D sky130_fd_sc_hd__or3_4
X_12645_ _12587_/Y _12607_/Y _12644_/X VGND VGND VPWR VPWR _12700_/A sky130_fd_sc_hd__or3_4
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24081__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11512__A _23759_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15364_ _15363_/Y _15359_/X _11576_/X _15359_/X VGND VGND VPWR VPWR _15364_/X sky130_fd_sc_hd__a2bb2o_4
X_18152_ _18152_/A VGND VGND VPWR VPWR _18316_/A sky130_fd_sc_hd__inv_2
XANTENNA__21846__B1 _24550_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12576_ _25044_/Q _24509_/Q _12647_/C _12575_/Y VGND VGND VPWR VPWR _12576_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20825__A _21097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24010__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14315_ _20177_/A _24780_/Q _14315_/C VGND VGND VPWR VPWR _14317_/B sky130_fd_sc_hd__or3_4
X_17103_ _17102_/X VGND VGND VPWR VPWR _17103_/Y sky130_fd_sc_hd__inv_2
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11527_ _11500_/X VGND VGND VPWR VPWR _11527_/Y sky130_fd_sc_hd__inv_2
X_18083_ _11733_/B _18080_/A VGND VGND VPWR VPWR _18086_/A sky130_fd_sc_hd__and2_4
XFILLER_129_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15919__A _15655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15525__B1 _14304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15295_ _15295_/A _15294_/Y VGND VGND VPWR VPWR _23761_/D sky130_fd_sc_hd__nor2_4
X_17034_ _17034_/A _17145_/A _17034_/C _17033_/X VGND VGND VPWR VPWR _17034_/X sky130_fd_sc_hd__or4_4
X_14246_ _14009_/Y _14243_/X _14218_/X _14226_/A VGND VGND VPWR VPWR _14246_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19806__A3 _15704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14542__B _14482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21074__B2 _11529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14177_ MSO_S3 _14176_/X _24830_/Q _14171_/X VGND VGND VPWR VPWR _14177_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__25216__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13128_ _13166_/A _23596_/Q VGND VGND VPWR VPWR _13128_/X sky130_fd_sc_hd__or2_4
XFILLER_3_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18985_ _18984_/Y _18982_/X _18938_/X _18982_/X VGND VGND VPWR VPWR _18985_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15654__A _15653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13059_ _11732_/A VGND VGND VPWR VPWR _13238_/A sky130_fd_sc_hd__buf_2
X_17936_ _17968_/A _17936_/B _17936_/C VGND VGND VPWR VPWR _17936_/X sky130_fd_sc_hd__and3_4
XFILLER_6_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17867_ _17899_/A _23530_/Q VGND VGND VPWR VPWR _17869_/B sky130_fd_sc_hd__or2_4
XFILLER_94_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19606_ _19606_/A VGND VGND VPWR VPWR _19606_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13174__A _13136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16818_ _16920_/A VGND VGND VPWR VPWR _16879_/A sky130_fd_sc_hd__buf_2
X_17798_ _17961_/A _17795_/X _17798_/C VGND VGND VPWR VPWR _17798_/X sky130_fd_sc_hd__and3_4
XFILLER_19_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24851__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19537_ _19536_/Y _19534_/X _11839_/X _19534_/X VGND VGND VPWR VPWR _23301_/D sky130_fd_sc_hd__a2bb2o_4
X_16749_ _24392_/Q VGND VGND VPWR VPWR _16749_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14802__A2_N _24126_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24169__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20888__B2 _11527_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19468_ _19467_/Y VGND VGND VPWR VPWR _19468_/X sky130_fd_sc_hd__buf_2
XFILLER_59_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18419_ _18419_/A VGND VGND VPWR VPWR _18427_/A sky130_fd_sc_hd__inv_2
X_19399_ _13106_/B VGND VGND VPWR VPWR _19399_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22934__B _22870_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21430_ _24030_/Q _20818_/X VGND VGND VPWR VPWR _21430_/X sky130_fd_sc_hd__or2_4
XANTENNA__21837__B1 _20782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21301__A2 _20931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22922__A1_N _12401_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21361_ _20892_/X _21359_/X _18011_/A _22548_/A VGND VGND VPWR VPWR _21361_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15516__B1 _15386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23100_ _23100_/CLK _20080_/X VGND VGND VPWR VPWR _23100_/Q sky130_fd_sc_hd__dfxtp_4
X_20312_ _14259_/Y _20296_/X _20286_/X _20311_/X VGND VGND VPWR VPWR _20313_/A sky130_fd_sc_hd__a211o_4
X_24080_ _24079_/CLK _24080_/D HRESETn VGND VGND VPWR VPWR _16760_/A sky130_fd_sc_hd__dfrtp_4
X_21292_ _21292_/A VGND VGND VPWR VPWR _21292_/X sky130_fd_sc_hd__buf_2
XFILLER_116_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23733__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23031_ _23011_/X _23015_/X _23030_/X VGND VGND VPWR VPWR HRDATA[31] sky130_fd_sc_hd__a21o_4
X_20243_ _13800_/A _20240_/X _20243_/C VGND VGND VPWR VPWR _20243_/X sky130_fd_sc_hd__or3_4
XFILLER_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20174_ _13891_/A _20161_/X _20165_/Y _20173_/X VGND VGND VPWR VPWR _20251_/B sky130_fd_sc_hd__a211o_4
XFILLER_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12084__A2_N _24561_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24982_ _24984_/CLK _24982_/D HRESETn VGND VGND VPWR VPWR _13370_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_131_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24939__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23933_ _24735_/CLK _23933_/D HRESETn VGND VGND VPWR VPWR _23933_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13084__A _13169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23864_ _23859_/CLK _23864_/D HRESETn VGND VGND VPWR VPWR _23864_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24592__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22815_ _22195_/X _22814_/X _22629_/X _24570_/Q _22198_/X VGND VGND VPWR VPWR _22816_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16395__A _16401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22868__A2 _22285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23795_ _23796_/CLK _20695_/X HRESETn VGND VGND VPWR VPWR _23795_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19194__B1 _19149_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24521__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23005__B _22015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22746_ _24278_/Q _22616_/X _22338_/X VGND VGND VPWR VPWR _22746_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14942__A1_N _14941_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15755__B1 _15332_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22677_ _22677_/A _22674_/X _22676_/X VGND VGND VPWR VPWR _22686_/A sky130_fd_sc_hd__and3_4
XFILLER_90_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22844__B _22015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12430_ _12418_/C _12417_/B _12401_/B _12417_/A VGND VGND VPWR VPWR _12433_/B sky130_fd_sc_hd__or4_4
X_24416_ _24425_/CLK _15856_/X HRESETn VGND VGND VPWR VPWR _24416_/Q sky130_fd_sc_hd__dfrtp_4
X_21628_ _21612_/A _19696_/Y VGND VGND VPWR VPWR _21630_/B sky130_fd_sc_hd__or2_4
X_12361_ _12495_/A _22373_/A _12360_/A _22373_/A VGND VGND VPWR VPWR _12361_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24347_ _23872_/CLK _16067_/X HRESETn VGND VGND VPWR VPWR _24347_/Q sky130_fd_sc_hd__dfrtp_4
X_21559_ _21308_/X _21552_/X _21080_/Y _21558_/X VGND VGND VPWR VPWR _21559_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_126_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14100_ _15260_/A VGND VGND VPWR VPWR _14100_/X sky130_fd_sc_hd__buf_2
X_15080_ _15059_/X VGND VGND VPWR VPWR _15080_/Y sky130_fd_sc_hd__inv_2
X_12292_ _12265_/B _12300_/A VGND VGND VPWR VPWR _12293_/B sky130_fd_sc_hd__or2_4
XFILLER_14_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16180__B1 _16179_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19249__B2 _19244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24278_ _24104_/CLK _16253_/X HRESETn VGND VGND VPWR VPWR _24278_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14031_ _20239_/A _14026_/X _13665_/X _14028_/X VGND VGND VPWR VPWR _14031_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17954__A _17725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14730__A1 _24706_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23229_ _23293_/CLK _19741_/X VGND VGND VPWR VPWR _19740_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__14730__B2 _14729_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20803__A1 _24500_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20803__B2 _15642_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17680__B1 _16678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22005__B1 _14732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18770_ _18768_/Y _18762_/X _18744_/X _18769_/X VGND VGND VPWR VPWR _18770_/X sky130_fd_sc_hd__a2bb2o_4
X_15982_ HWDATA[8] VGND VGND VPWR VPWR _15982_/X sky130_fd_sc_hd__buf_2
XANTENNA__21359__A2 _14016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17721_ _17721_/A VGND VGND VPWR VPWR _17881_/A sky130_fd_sc_hd__buf_2
X_14933_ _24272_/Q VGND VGND VPWR VPWR _14933_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24609__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17652_ _21335_/A _17626_/X _17648_/X VGND VGND VPWR VPWR _17652_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_8_113_0_HCLK clkbuf_7_56_0_HCLK/X VGND VGND VPWR VPWR _23676_/CLK sky130_fd_sc_hd__clkbuf_1
X_14864_ _14693_/Y _15016_/A _14830_/X _14863_/X VGND VGND VPWR VPWR _14864_/X sky130_fd_sc_hd__o22a_4
XFILLER_91_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14246__B1 _14218_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16603_ _16601_/Y _16595_/X _15507_/X _16602_/X VGND VGND VPWR VPWR _16603_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_176_0_HCLK clkbuf_7_88_0_HCLK/X VGND VGND VPWR VPWR _24523_/CLK sky130_fd_sc_hd__clkbuf_1
X_13815_ _13815_/A VGND VGND VPWR VPWR _13815_/X sky130_fd_sc_hd__buf_2
X_14795_ _14750_/X _14794_/X VGND VGND VPWR VPWR _14982_/A sky130_fd_sc_hd__or2_4
X_17583_ _17494_/Y _17577_/X _17528_/X _17580_/B VGND VGND VPWR VPWR _17583_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15994__B1 _15992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22100__A _20961_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14818__A _14818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24262__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19185__B1 _19095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19322_ _19321_/Y _19319_/X _19207_/X _19319_/X VGND VGND VPWR VPWR _23376_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13746_ _13716_/A VGND VGND VPWR VPWR _13769_/A sky130_fd_sc_hd__buf_2
X_16534_ _16534_/A VGND VGND VPWR VPWR _16534_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22457__D _22456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21531__A2 _14016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19253_ _23400_/Q VGND VGND VPWR VPWR _21169_/B sky130_fd_sc_hd__inv_2
X_13677_ _20201_/A _20201_/B _13677_/C VGND VGND VPWR VPWR _13677_/X sky130_fd_sc_hd__or3_4
X_16465_ _16401_/A VGND VGND VPWR VPWR _16465_/X sky130_fd_sc_hd__buf_2
XANTENNA__24770__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18204_ _23859_/Q VGND VGND VPWR VPWR _18205_/D sky130_fd_sc_hd__inv_2
X_12628_ _25043_/Q VGND VGND VPWR VPWR _12739_/A sky130_fd_sc_hd__inv_2
X_15416_ _13644_/A VGND VGND VPWR VPWR _15416_/X sky130_fd_sc_hd__buf_2
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16396_ _16395_/X VGND VGND VPWR VPWR _16396_/X sky130_fd_sc_hd__buf_2
X_19184_ _23424_/Q VGND VGND VPWR VPWR _19184_/Y sky130_fd_sc_hd__inv_2
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21295__A1 _24397_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15347_ _15347_/A VGND VGND VPWR VPWR _15347_/Y sky130_fd_sc_hd__inv_2
X_18135_ _16111_/A _18318_/A _16056_/Y _18244_/A VGND VGND VPWR VPWR _18135_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12792__A1_N _22712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12559_ _24523_/Q VGND VGND VPWR VPWR _12559_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22492__B1 _16649_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18160__A1 _16121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15278_ _24629_/Q VGND VGND VPWR VPWR _15278_/Y sky130_fd_sc_hd__inv_2
X_18066_ _19801_/B VGND VGND VPWR VPWR _18067_/A sky130_fd_sc_hd__buf_2
XFILLER_117_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16171__B1 _15772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14229_ _14223_/Y _14226_/X _14228_/X _14226_/X VGND VGND VPWR VPWR _14229_/X sky130_fd_sc_hd__a2bb2o_4
X_17017_ _17017_/A _17017_/B _17017_/C _17016_/X VGND VGND VPWR VPWR _17017_/X sky130_fd_sc_hd__or4_4
XANTENNA__13169__A _13169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25050__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22795__A1 _15846_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22795__B2 _21543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21386__A _21229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18968_ _18968_/A _18072_/X _20134_/C VGND VGND VPWR VPWR _18969_/A sky130_fd_sc_hd__or3_4
XFILLER_113_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17919_ _17887_/A _19206_/A VGND VGND VPWR VPWR _17921_/B sky130_fd_sc_hd__or2_4
X_18899_ _18898_/X VGND VGND VPWR VPWR _18899_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_72_0_HCLK clkbuf_7_73_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_72_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20930_ _20910_/X _20925_/Y _20927_/X _20929_/X VGND VGND VPWR VPWR _20930_/X sky130_fd_sc_hd__a211o_4
XFILLER_94_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20861_ _15159_/A _20861_/B VGND VGND VPWR VPWR _20861_/X sky130_fd_sc_hd__and2_4
XANTENNA__15985__B1 _15890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14788__B2 _24123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22010__A _21886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19176__B1 _19152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14728__A _24706_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22600_ _22599_/X VGND VGND VPWR VPWR _22600_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23580_ _23563_/CLK _23580_/D VGND VGND VPWR VPWR _18742_/A sky130_fd_sc_hd__dfxtp_4
X_20792_ _20759_/X _20791_/X _20737_/B _12062_/X VGND VGND VPWR VPWR _20792_/X sky130_fd_sc_hd__o22a_4
XPHY_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18923__B1 _18901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22531_ _21069_/X VGND VGND VPWR VPWR _22531_/X sky130_fd_sc_hd__buf_2
XFILLER_23_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14756__A2_N _14754_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21315__A2_N _14015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23985__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22462_ _22256_/B _22461_/X VGND VGND VPWR VPWR _22462_/X sky130_fd_sc_hd__and2_4
XFILLER_50_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20465__A _20465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24201_ _24201_/CLK _24201_/D HRESETn VGND VGND VPWR VPWR _24201_/Q sky130_fd_sc_hd__dfrtp_4
X_21413_ _21413_/A VGND VGND VPWR VPWR _21413_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23914__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15559__A _19455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25181_ _24847_/CLK _25181_/D HRESETn VGND VGND VPWR VPWR _17448_/B sky130_fd_sc_hd__dfrtp_4
X_22393_ _20748_/X _22390_/Y _21029_/X _22392_/X VGND VGND VPWR VPWR _22394_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25138__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24132_ _24098_/CLK _16609_/X HRESETn VGND VGND VPWR VPWR _16608_/A sky130_fd_sc_hd__dfrtp_4
X_21344_ _21158_/A _21344_/B VGND VGND VPWR VPWR _21344_/X sky130_fd_sc_hd__or2_4
XFILLER_136_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24063_ _24064_/CLK _16946_/Y HRESETn VGND VGND VPWR VPWR _16835_/A sky130_fd_sc_hd__dfrtp_4
X_21275_ _21275_/A VGND VGND VPWR VPWR _21276_/A sky130_fd_sc_hd__inv_2
XFILLER_11_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22786__A1 _12448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11526__B2 _11521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21589__A2 _22840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22786__B2 _20747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23014_ _12305_/Y _22259_/X _24058_/Q _22433_/A VGND VGND VPWR VPWR _23015_/D sky130_fd_sc_hd__a2bb2o_4
X_20226_ _14012_/Y _20217_/Y _20254_/A VGND VGND VPWR VPWR _20226_/X sky130_fd_sc_hd__and3_4
XFILLER_81_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22830__D _22829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21296__A _22167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15610__A1_N _12592_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20157_ _20156_/X VGND VGND VPWR VPWR _20157_/X sky130_fd_sc_hd__buf_2
XFILLER_89_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24773__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22538__B2 _22537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24965_ _24980_/CLK _24965_/D HRESETn VGND VGND VPWR VPWR _24965_/Q sky130_fd_sc_hd__dfrtp_4
X_20088_ _20088_/A VGND VGND VPWR VPWR _21332_/B sky130_fd_sc_hd__inv_2
XANTENNA__24702__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11930_ _11930_/A VGND VGND VPWR VPWR _11930_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23916_ _24928_/CLK _23916_/D HRESETn VGND VGND VPWR VPWR _21871_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24896_ _24902_/CLK _13920_/X HRESETn VGND VGND VPWR VPWR _13815_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_17_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11861_ _11859_/Y _11852_/X _11860_/X _11830_/Y VGND VGND VPWR VPWR _25169_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15741__B _15741_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23016__A _24124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23847_ _23845_/CLK _23847_/D HRESETn VGND VGND VPWR VPWR _18159_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15976__B1 _15788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_249_0_HCLK clkbuf_7_124_0_HCLK/X VGND VGND VPWR VPWR _24113_/CLK sky130_fd_sc_hd__clkbuf_1
X_13600_ _11663_/Y _13555_/X VGND VGND VPWR VPWR _13600_/Y sky130_fd_sc_hd__nand2_4
X_14580_ _17698_/A _14561_/A _14573_/X VGND VGND VPWR VPWR _24735_/D sky130_fd_sc_hd__a21oi_4
X_11792_ _25184_/Q _11772_/B _11815_/C _11809_/B VGND VGND VPWR VPWR _11793_/A sky130_fd_sc_hd__a211o_4
XFILLER_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23778_ _23668_/CLK _20187_/X HRESETn VGND VGND VPWR VPWR _20162_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_26_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13531_ _23732_/Q _13531_/B VGND VGND VPWR VPWR _13532_/B sky130_fd_sc_hd__or2_4
XFILLER_13_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22729_ _22547_/X _22727_/X _22551_/X _22728_/X VGND VGND VPWR VPWR _22730_/B sky130_fd_sc_hd__o22a_4
XFILLER_41_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22574__B _22574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16250_ _16228_/X _16234_/X _15596_/X _24280_/Q _16237_/X VGND VGND VPWR VPWR _16250_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_9_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13462_ _13462_/A _13461_/X VGND VGND VPWR VPWR _13463_/A sky130_fd_sc_hd__or2_4
XFILLER_90_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15201_ _15108_/B _15213_/B VGND VGND VPWR VPWR _15211_/B sky130_fd_sc_hd__or2_4
X_12413_ _12413_/A _12360_/A _12411_/X _12413_/D VGND VGND VPWR VPWR _12414_/B sky130_fd_sc_hd__or4_4
XANTENNA__21277__A1 _16121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11997__A _25144_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23655__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16181_ _16181_/A VGND VGND VPWR VPWR _16181_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13393_ _13392_/X VGND VGND VPWR VPWR _13393_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14951__B2 _22477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15132_ _15132_/A _15130_/A VGND VGND VPWR VPWR _15133_/C sky130_fd_sc_hd__or2_4
X_12344_ _12344_/A VGND VGND VPWR VPWR _12344_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23018__A2 _22505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15063_ _14694_/A _15063_/B VGND VGND VPWR VPWR _15063_/X sky130_fd_sc_hd__or2_4
X_19940_ _19938_/Y _19939_/X _15556_/X _19939_/X VGND VGND VPWR VPWR _19940_/X sky130_fd_sc_hd__a2bb2o_4
X_12275_ _12275_/A _12278_/B VGND VGND VPWR VPWR _12275_/Y sky130_fd_sc_hd__nand2_4
X_14014_ _15407_/A VGND VGND VPWR VPWR _14015_/A sky130_fd_sc_hd__buf_2
XFILLER_49_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20822__B _20821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19871_ _19871_/A VGND VGND VPWR VPWR _21683_/B sky130_fd_sc_hd__inv_2
XANTENNA__15916__B _15422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19642__B2 _19636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18822_ _18809_/A VGND VGND VPWR VPWR _18822_/X sky130_fd_sc_hd__buf_2
XFILLER_95_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22529__A1 _17498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14834__A1_N _15034_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18753_ _18751_/Y _18752_/X _18706_/X _18752_/X VGND VGND VPWR VPWR _23577_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15965_ _22436_/A VGND VGND VPWR VPWR _15965_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24443__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17704_ _17689_/X _17696_/X _17703_/X _15712_/X _15720_/X VGND VGND VPWR VPWR _17704_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_64_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_59_0_HCLK clkbuf_6_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_59_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14916_ _24262_/Q VGND VGND VPWR VPWR _14916_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18684_ _18684_/A VGND VGND VPWR VPWR _18684_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14219__B1 _14218_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21653__B _21653_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15896_ _24400_/Q VGND VGND VPWR VPWR _15896_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17635_ _23941_/Q VGND VGND VPWR VPWR _17636_/A sky130_fd_sc_hd__buf_2
X_14847_ _15019_/B _24137_/Q _15019_/B _24137_/Q VGND VGND VPWR VPWR _14847_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15967__B1 _11585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19158__B1 _19089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17566_ _16718_/A _17565_/Y VGND VGND VPWR VPWR _17566_/X sky130_fd_sc_hd__or2_4
X_14778_ _15059_/A _24097_/Q _24710_/Q _14777_/Y VGND VGND VPWR VPWR _14784_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14267__B _18633_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22701__A1 _22195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19305_ _19304_/Y VGND VGND VPWR VPWR _19305_/X sky130_fd_sc_hd__buf_2
XANTENNA__22701__B2 _22198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16517_ _24173_/Q VGND VGND VPWR VPWR _16517_/Y sky130_fd_sc_hd__inv_2
X_13729_ _13728_/X VGND VGND VPWR VPWR _13732_/B sky130_fd_sc_hd__inv_2
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17497_ _17497_/A _17497_/B _16692_/Y _17497_/D VGND VGND VPWR VPWR _17497_/X sky130_fd_sc_hd__or4_4
XANTENNA__22484__B _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19236_ _18030_/A _17625_/A _18022_/X VGND VGND VPWR VPWR _19236_/X sky130_fd_sc_hd__or3_4
XFILLER_32_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16448_ _16448_/A VGND VGND VPWR VPWR _16448_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19167_ _24732_/Q _19167_/B _19144_/A _19189_/B VGND VGND VPWR VPWR _19167_/X sky130_fd_sc_hd__or4_4
X_16379_ _16313_/A VGND VGND VPWR VPWR _16379_/X sky130_fd_sc_hd__buf_2
XANTENNA__14942__B2 _24269_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18118_ _18118_/A VGND VGND VPWR VPWR _18118_/X sky130_fd_sc_hd__buf_2
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19098_ _19097_/Y _19092_/X _18964_/X _19078_/Y VGND VGND VPWR VPWR _23455_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19881__B2 _19876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24628__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17594__A _16685_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18049_ _18048_/X VGND VGND VPWR VPWR _18049_/X sky130_fd_sc_hd__buf_2
XANTENNA__16695__B2 _20778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21060_ _13360_/A _21055_/X _21058_/X _24503_/Q _21059_/X VGND VGND VPWR VPWR _21060_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_67_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20011_ _23126_/Q _20010_/Y _23666_/D _20010_/A VGND VGND VPWR VPWR _23126_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13627__A _21448_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21440__B2 _21083_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12531__A _12534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16970__A1_N _24310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24184__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16938__A _16936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24750_ _24750_/CLK _24750_/D HRESETn VGND VGND VPWR VPWR _14511_/A sky130_fd_sc_hd__dfrtp_4
X_21962_ _21371_/A _21962_/B VGND VGND VPWR VPWR _21962_/X sky130_fd_sc_hd__or2_4
XFILLER_73_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24113__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22940__A1 _11524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23701_ _23702_/CLK _20445_/Y HRESETn VGND VGND VPWR VPWR _21887_/A sky130_fd_sc_hd__dfrtp_4
X_20913_ _19279_/A _14016_/A _19231_/A _20827_/X VGND VGND VPWR VPWR _20913_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22940__B2 _22537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15958__B1 _15777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24681_ _24681_/CLK _15122_/X HRESETn VGND VGND VPWR VPWR _24681_/Q sky130_fd_sc_hd__dfrtp_4
X_21893_ _11938_/A _21300_/B _24778_/Q _23622_/Q _22218_/C VGND VGND VPWR VPWR _21893_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_42_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13362__A _13362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23632_ _23641_/CLK _23632_/D HRESETn VGND VGND VPWR VPWR _20288_/A sky130_fd_sc_hd__dfrtp_4
X_20844_ _14064_/A _20844_/B VGND VGND VPWR VPWR _20849_/A sky130_fd_sc_hd__and2_4
XFILLER_74_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_2_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_16_0_HCLK clkbuf_7_8_0_HCLK/X VGND VGND VPWR VPWR _24847_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23563_ _23563_/CLK _23563_/D VGND VGND VPWR VPWR _18792_/A sky130_fd_sc_hd__dfxtp_4
X_20775_ _21850_/A VGND VGND VPWR VPWR _22438_/A sky130_fd_sc_hd__buf_2
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_79_0_HCLK clkbuf_8_79_0_HCLK/A VGND VGND VPWR VPWR _24776_/CLK sky130_fd_sc_hd__clkbuf_1
X_22514_ _21848_/B VGND VGND VPWR VPWR _22757_/B sky130_fd_sc_hd__buf_2
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23494_ _23493_/CLK _23494_/D VGND VGND VPWR VPWR _23494_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20195__A _20195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22445_ _24139_/Q _22445_/B VGND VGND VPWR VPWR _22445_/X sky130_fd_sc_hd__and2_4
XANTENNA__14193__A _20195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12944__B1 _12896_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11610__A _11599_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25164_ _24623_/CLK _25164_/D HRESETn VGND VGND VPWR VPWR _11879_/A sky130_fd_sc_hd__dfrtp_4
X_22376_ _22376_/A _21850_/A VGND VGND VPWR VPWR _22379_/B sky130_fd_sc_hd__and2_4
XFILLER_135_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22208__B1 _16450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24115_ _24698_/CLK _24115_/D HRESETn VGND VGND VPWR VPWR _24115_/Q sky130_fd_sc_hd__dfrtp_4
X_21327_ _21130_/X _21325_/X _21326_/X VGND VGND VPWR VPWR _21327_/X sky130_fd_sc_hd__and3_4
XANTENNA__16686__B2 _16693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25095_ _25097_/CLK _25095_/D HRESETn VGND VGND VPWR VPWR _25095_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24954__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12060_ _12060_/A VGND VGND VPWR VPWR _12061_/B sky130_fd_sc_hd__buf_2
X_24046_ _24308_/CLK _17106_/X HRESETn VGND VGND VPWR VPWR _24046_/Q sky130_fd_sc_hd__dfrtp_4
X_21258_ _22146_/B _21255_/X _21256_/X _21257_/X VGND VGND VPWR VPWR _21259_/A sky130_fd_sc_hd__a211o_4
XFILLER_81_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15736__B _16127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20209_ _20209_/A _20209_/B VGND VGND VPWR VPWR _20209_/X sky130_fd_sc_hd__or2_4
XFILLER_137_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21189_ _22806_/B _21185_/X _20745_/X _21188_/X VGND VGND VPWR VPWR _21189_/X sky130_fd_sc_hd__a211o_4
XANTENNA__12441__A _12434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19388__B1 _19387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12962_ _12867_/X VGND VGND VPWR VPWR _12992_/A sky130_fd_sc_hd__buf_2
X_15750_ _15744_/X VGND VGND VPWR VPWR _15750_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24948_ _23925_/CLK _24948_/D HRESETn VGND VGND VPWR VPWR _11676_/A sky130_fd_sc_hd__dfrtp_4
X_11913_ _24986_/Q VGND VGND VPWR VPWR _11913_/Y sky130_fd_sc_hd__inv_2
X_14701_ _24688_/Q _14699_/Y _14881_/A _14714_/A VGND VGND VPWR VPWR _14705_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12893_ _12886_/X _12892_/X VGND VGND VPWR VPWR _12894_/B sky130_fd_sc_hd__or2_4
X_15681_ _12339_/Y _15677_/X _11566_/X _15680_/X VGND VGND VPWR VPWR _24486_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15949__B1 _15855_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24879_ _24879_/CLK _14029_/X HRESETn VGND VGND VPWR VPWR _20232_/A sky130_fd_sc_hd__dfrtp_4
X_17420_ _17262_/Y _17423_/B VGND VGND VPWR VPWR _17420_/Y sky130_fd_sc_hd__nand2_4
X_11844_ _19603_/A VGND VGND VPWR VPWR _11844_/X sky130_fd_sc_hd__buf_2
X_14632_ _15270_/A _14621_/X _14622_/X _14631_/Y VGND VGND VPWR VPWR _14632_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23836__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14563_ _14563_/A VGND VGND VPWR VPWR _17947_/A sky130_fd_sc_hd__buf_2
X_17351_ _17353_/B VGND VGND VPWR VPWR _17352_/B sky130_fd_sc_hd__inv_2
X_11775_ _11771_/Y _11694_/X VGND VGND VPWR VPWR _11802_/C sky130_fd_sc_hd__or2_4
XFILLER_57_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16302_ _16302_/A _16306_/B VGND VGND VPWR VPWR _16302_/Y sky130_fd_sc_hd__nor2_4
XFILLER_9_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13514_ _13513_/X VGND VGND VPWR VPWR _13514_/X sky130_fd_sc_hd__buf_2
XFILLER_105_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14494_ _14469_/X VGND VGND VPWR VPWR _14494_/X sky130_fd_sc_hd__buf_2
X_17282_ _17278_/X _17279_/X _17280_/X _17282_/D VGND VGND VPWR VPWR _17296_/B sky130_fd_sc_hd__or4_4
XANTENNA__16374__B1 _16373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19021_ _21663_/B _19018_/X _15554_/X _19018_/X VGND VGND VPWR VPWR _19021_/X sky130_fd_sc_hd__a2bb2o_4
X_13445_ _22483_/A _24768_/Q _22483_/A _24768_/Q VGND VGND VPWR VPWR _13453_/B sky130_fd_sc_hd__a2bb2o_4
X_16233_ _16625_/A VGND VGND VPWR VPWR _16234_/A sky130_fd_sc_hd__buf_2
XFILLER_103_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11520__A _11599_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13376_ _13376_/A VGND VGND VPWR VPWR _13376_/Y sky130_fd_sc_hd__inv_2
X_16164_ _24310_/Q VGND VGND VPWR VPWR _16164_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16126__B1 _15291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20833__A _22858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12327_ _25088_/Q _22591_/A _12412_/A _12326_/Y VGND VGND VPWR VPWR _12327_/X sky130_fd_sc_hd__o22a_4
X_15115_ _15115_/A _15159_/B VGND VGND VPWR VPWR _15115_/X sky130_fd_sc_hd__or2_4
X_16095_ _24336_/Q VGND VGND VPWR VPWR _16095_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24695__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15046_ _15018_/X _15046_/B _15046_/C VGND VGND VPWR VPWR _15046_/X sky130_fd_sc_hd__and3_4
X_19923_ _19922_/Y _19918_/X _19859_/X _19918_/A VGND VGND VPWR VPWR _19923_/X sky130_fd_sc_hd__a2bb2o_4
X_12258_ _12257_/X VGND VGND VPWR VPWR _12259_/B sky130_fd_sc_hd__inv_2
XFILLER_64_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24624__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19854_ _19841_/X VGND VGND VPWR VPWR _19854_/X sky130_fd_sc_hd__buf_2
XFILLER_25_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12189_ _12073_/Y _12189_/B VGND VGND VPWR VPWR _12190_/C sky130_fd_sc_hd__or2_4
X_18805_ _18804_/Y _18798_/X _18712_/X _18798_/A VGND VGND VPWR VPWR _23559_/D sky130_fd_sc_hd__a2bb2o_4
X_19785_ _23212_/Q VGND VGND VPWR VPWR _21778_/B sky130_fd_sc_hd__inv_2
X_16997_ _16188_/Y _24039_/Q _16188_/Y _24039_/Q VGND VGND VPWR VPWR _16997_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19379__B1 _19311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22479__B _22265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18736_ _18752_/A VGND VGND VPWR VPWR _18736_/X sky130_fd_sc_hd__buf_2
XFILLER_114_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15948_ _15928_/X VGND VGND VPWR VPWR _15948_/X sky130_fd_sc_hd__buf_2
XFILLER_23_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18667_ _18666_/X VGND VGND VPWR VPWR _18682_/A sky130_fd_sc_hd__inv_2
X_15879_ _24406_/Q VGND VGND VPWR VPWR _15879_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13182__A _13182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17618_ _17615_/A _17615_/B VGND VGND VPWR VPWR _17618_/Y sky130_fd_sc_hd__nand2_4
X_18598_ _16358_/Y _18338_/X _16378_/A _18427_/A VGND VGND VPWR VPWR _18598_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_232_0_HCLK clkbuf_8_233_0_HCLK/A VGND VGND VPWR VPWR _25090_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17549_ _17497_/A _17497_/B _17548_/X VGND VGND VPWR VPWR _17550_/B sky130_fd_sc_hd__or3_4
XANTENNA__16493__A _16493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20560_ _16553_/Y _20553_/X _20556_/X _20559_/Y VGND VGND VPWR VPWR _20560_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16365__B1 _15978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15707__A3 _15706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19219_ _21746_/A _19213_/X _19152_/X _19218_/X VGND VGND VPWR VPWR _19219_/X sky130_fd_sc_hd__a2bb2o_4
X_20491_ _20499_/C _20517_/A VGND VGND VPWR VPWR _20491_/X sky130_fd_sc_hd__or2_4
X_22230_ _22230_/A VGND VGND VPWR VPWR _22551_/A sky130_fd_sc_hd__buf_2
XFILLER_69_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21839__A _21839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20743__A _21113_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22161_ _22161_/A _22953_/B VGND VGND VPWR VPWR _22161_/X sky130_fd_sc_hd__and2_4
XANTENNA__15837__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14679__B1 _24867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21112_ _20926_/A _21109_/X _22279_/A _21111_/X VGND VGND VPWR VPWR _21112_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14143__A2 _13492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22092_ _21617_/A _22092_/B VGND VGND VPWR VPWR _22092_/X sky130_fd_sc_hd__or2_4
XFILLER_87_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24365__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21043_ _22036_/A VGND VGND VPWR VPWR _21043_/X sky130_fd_sc_hd__buf_2
XANTENNA__13357__A _11503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13367__A1_N _22006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15572__A _15572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24802_ _24811_/CLK _24802_/D HRESETn VGND VGND VPWR VPWR _14259_/A sky130_fd_sc_hd__dfstp_4
XFILLER_41_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22994_ _21864_/X _22992_/X _22530_/X _22993_/X VGND VGND VPWR VPWR _22994_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14851__B1 _24706_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_42_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_42_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21945_ _21941_/X _21944_/X _14488_/X VGND VGND VPWR VPWR _21945_/Y sky130_fd_sc_hd__o21ai_4
X_24733_ _24733_/CLK _24733_/D HRESETn VGND VGND VPWR VPWR _24733_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18883__A _18743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13092__A _13092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24664_ _24671_/CLK _24664_/D HRESETn VGND VGND VPWR VPWR _24664_/Q sky130_fd_sc_hd__dfrtp_4
X_21876_ _21876_/A _15639_/X VGND VGND VPWR VPWR _21876_/X sky130_fd_sc_hd__and2_4
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23615_ _24013_/CLK _20269_/X HRESETn VGND VGND VPWR VPWR _23615_/Q sky130_fd_sc_hd__dfrtp_4
X_20827_ _15637_/X VGND VGND VPWR VPWR _20827_/X sky130_fd_sc_hd__buf_2
XPHY_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25153__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24595_ _24596_/CLK _24595_/D HRESETn VGND VGND VPWR VPWR _24595_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ _11557_/Y _11551_/X _11558_/X _11559_/X VGND VGND VPWR VPWR _25212_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_51_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23546_ _23479_/CLK _18843_/X VGND VGND VPWR VPWR _23546_/Q sky130_fd_sc_hd__dfxtp_4
X_20758_ _20861_/B VGND VGND VPWR VPWR _20758_/X sky130_fd_sc_hd__buf_2
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23477_ _23537_/CLK _23477_/D VGND VGND VPWR VPWR _13097_/B sky130_fd_sc_hd__dfxtp_4
X_20689_ _11900_/A _20691_/B VGND VGND VPWR VPWR _23786_/D sky130_fd_sc_hd__and2_4
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _13230_/A _23129_/Q VGND VGND VPWR VPWR _13231_/C sky130_fd_sc_hd__or2_4
XFILLER_109_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25216_ _24385_/CLK _11546_/X HRESETn VGND VGND VPWR VPWR _25216_/Q sky130_fd_sc_hd__dfrtp_4
X_22428_ _21434_/A VGND VGND VPWR VPWR _22433_/A sky130_fd_sc_hd__buf_2
XANTENNA__16108__B1 _15982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21101__B1 _22858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13161_ _13261_/A _13161_/B VGND VGND VPWR VPWR _13161_/X sky130_fd_sc_hd__or2_4
XANTENNA__21652__A1 _22745_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12393__B2 _21567_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25147_ _24984_/CLK _25147_/D HRESETn VGND VGND VPWR VPWR _25147_/Q sky130_fd_sc_hd__dfrtp_4
X_22359_ _22348_/X _22349_/X _22353_/X _22354_/Y _22358_/Y VGND VGND VPWR VPWR _22381_/C
+ sky130_fd_sc_hd__a32o_4
XFILLER_136_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12112_ _12110_/A _24554_/Q _12176_/A _12111_/Y VGND VGND VPWR VPWR _12119_/B sky130_fd_sc_hd__o22a_4
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13092_ _13092_/A _23373_/Q VGND VGND VPWR VPWR _13092_/X sky130_fd_sc_hd__or2_4
X_25078_ _25090_/CLK _12519_/X HRESETn VGND VGND VPWR VPWR _12328_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_123_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13342__B1 _11616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12043_ _12039_/A _12035_/X _12041_/Y VGND VGND VPWR VPWR _12043_/X sky130_fd_sc_hd__o21a_4
X_16920_ _16920_/A _16837_/D VGND VGND VPWR VPWR _16921_/D sky130_fd_sc_hd__or2_4
XANTENNA__13267__A _13299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21404__A1 _22146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24029_ _24590_/CLK _24029_/D HRESETn VGND VGND VPWR VPWR _21291_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24035__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_124_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_124_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_16851_ _16850_/X VGND VGND VPWR VPWR _24089_/D sky130_fd_sc_hd__inv_2
XFILLER_38_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15802_ _12819_/Y _15795_/X _15801_/X _15757_/A VGND VGND VPWR VPWR _15802_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15482__A _11532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19570_ _21158_/B _19567_/X _11860_/X _19567_/X VGND VGND VPWR VPWR _23288_/D sky130_fd_sc_hd__a2bb2o_4
X_16782_ _16775_/X _16782_/B _16782_/C _16781_/X VGND VGND VPWR VPWR _16783_/D sky130_fd_sc_hd__or4_4
X_13994_ _13993_/X VGND VGND VPWR VPWR _13994_/Y sky130_fd_sc_hd__inv_2
X_18521_ _18520_/X VGND VGND VPWR VPWR _23825_/D sky130_fd_sc_hd__inv_2
XFILLER_74_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15733_ _13474_/B _15729_/X VGND VGND VPWR VPWR _15733_/X sky130_fd_sc_hd__and2_4
X_12945_ _12809_/Y _12943_/X _12944_/Y VGND VGND VPWR VPWR _25024_/D sky130_fd_sc_hd__o21a_4
XFILLER_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11515__A _11514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18452_ _18459_/A _18438_/X _18452_/C _18462_/A VGND VGND VPWR VPWR _18453_/A sky130_fd_sc_hd__or4_4
X_15664_ _15664_/A VGND VGND VPWR VPWR _15695_/A sky130_fd_sc_hd__inv_2
XANTENNA__21931__B _21931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12876_ _12876_/A _12805_/Y VGND VGND VPWR VPWR _12876_/X sky130_fd_sc_hd__or2_4
X_17403_ _17315_/Y _17400_/X VGND VGND VPWR VPWR _17404_/C sky130_fd_sc_hd__or2_4
XANTENNA__23670__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14615_ _14615_/A VGND VGND VPWR VPWR _14615_/Y sky130_fd_sc_hd__inv_2
X_11827_ _19597_/A VGND VGND VPWR VPWR _11827_/Y sky130_fd_sc_hd__inv_2
X_18383_ _16471_/A _18551_/A _16462_/A _18421_/B VGND VGND VPWR VPWR _18383_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22668__B1 _13362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15595_ _15574_/X _15582_/X _15477_/X _24528_/Q _15585_/X VGND VGND VPWR VPWR _15595_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17362_/A _17332_/X _17334_/C VGND VGND VPWR VPWR _24009_/D sky130_fd_sc_hd__and3_4
XANTENNA__17202__A _16373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11755_/Y _18075_/A _17227_/B VGND VGND VPWR VPWR _11758_/X sky130_fd_sc_hd__a21o_4
X_14546_ _14541_/D VGND VGND VPWR VPWR _19883_/B sky130_fd_sc_hd__buf_2
XFILLER_81_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_62_0_HCLK clkbuf_8_63_0_HCLK/A VGND VGND VPWR VPWR _24378_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17265_ _25192_/Q _17264_/A _11633_/Y _17264_/Y VGND VGND VPWR VPWR _17265_/X sky130_fd_sc_hd__o22a_4
X_11689_ _11687_/A _23912_/Q _11687_/Y _11688_/Y VGND VGND VPWR VPWR _11689_/X sky130_fd_sc_hd__o22a_4
X_14477_ _14437_/A VGND VGND VPWR VPWR _14482_/A sky130_fd_sc_hd__inv_2
XANTENNA__12346__A _12346_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19004_ _19002_/Y _19003_/X _15563_/X _19003_/X VGND VGND VPWR VPWR _19004_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24876__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16216_ _16216_/A VGND VGND VPWR VPWR _16216_/X sky130_fd_sc_hd__buf_2
X_13428_ _13428_/A VGND VGND VPWR VPWR _13428_/Y sky130_fd_sc_hd__inv_2
X_17196_ _14618_/A VGND VGND VPWR VPWR _20401_/A sky130_fd_sc_hd__buf_2
XFILLER_31_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13359_ _13358_/X VGND VGND VPWR VPWR _13360_/A sky130_fd_sc_hd__buf_2
X_16147_ _24317_/Q VGND VGND VPWR VPWR _16147_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21643__B2 _21181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21271__A1_N _21040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16078_ _16078_/A VGND VGND VPWR VPWR _16078_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15029_ _15029_/A VGND VGND VPWR VPWR _15029_/Y sky130_fd_sc_hd__inv_2
X_19906_ _19918_/A VGND VGND VPWR VPWR _19906_/X sky130_fd_sc_hd__buf_2
XFILLER_69_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19837_ _23191_/Q VGND VGND VPWR VPWR _19837_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21394__A _21394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19768_ _21609_/B _19765_/X _19721_/X _19765_/X VGND VGND VPWR VPWR _19768_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18719_ _18719_/A VGND VGND VPWR VPWR _18719_/X sky130_fd_sc_hd__buf_2
XANTENNA__23758__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_29_0_HCLK clkbuf_4_14_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19699_ _19698_/Y _19694_/X _19610_/X _19694_/X VGND VGND VPWR VPWR _23242_/D sky130_fd_sc_hd__a2bb2o_4
X_21730_ _21562_/A _21728_/X _21280_/X _21729_/X VGND VGND VPWR VPWR _21730_/X sky130_fd_sc_hd__o22a_4
XFILLER_24_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16586__B1 _16334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21661_ _21656_/X _21660_/X _14486_/X VGND VGND VPWR VPWR _21672_/B sky130_fd_sc_hd__o21a_4
XFILLER_71_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23400_ _23385_/CLK _23400_/D VGND VGND VPWR VPWR _23400_/Q sky130_fd_sc_hd__dfxtp_4
X_20612_ _20609_/Y _20610_/Y _20611_/X VGND VGND VPWR VPWR _20612_/X sky130_fd_sc_hd__o21a_4
X_24380_ _24378_/CLK _24380_/D HRESETn VGND VGND VPWR VPWR _24380_/Q sky130_fd_sc_hd__dfrtp_4
X_21592_ _21298_/B _21592_/B _21591_/X VGND VGND VPWR VPWR _21592_/X sky130_fd_sc_hd__and3_4
XANTENNA__21331__B1 _18049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23331_ _23313_/CLK _23331_/D VGND VGND VPWR VPWR _19451_/A sky130_fd_sc_hd__dfxtp_4
X_20543_ _20541_/Y _20538_/Y _20542_/X VGND VGND VPWR VPWR _20543_/X sky130_fd_sc_hd__o21a_4
XFILLER_137_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15010__B1 _14984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12375__A2_N _24482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21569__A _21569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23262_ _23278_/CLK _19648_/X VGND VGND VPWR VPWR _19643_/A sky130_fd_sc_hd__dfxtp_4
X_20474_ _13508_/D _20469_/X VGND VGND VPWR VPWR _20474_/X sky130_fd_sc_hd__or2_4
XFILLER_10_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24546__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25001_ _24998_/CLK _25001_/D HRESETn VGND VGND VPWR VPWR _25001_/Q sky130_fd_sc_hd__dfrtp_4
X_22213_ _21870_/A _22211_/X _21886_/X _22212_/X VGND VGND VPWR VPWR _22213_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12375__B2 _24482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23193_ _25106_/CLK _19833_/X VGND VGND VPWR VPWR _23193_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22144_ _22144_/A VGND VGND VPWR VPWR _22183_/A sky130_fd_sc_hd__inv_2
XFILLER_106_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22075_ _22055_/X _22075_/B VGND VGND VPWR VPWR _22075_/X sky130_fd_sc_hd__or2_4
XFILLER_121_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21026_ _20908_/X _20920_/X _20930_/X _20939_/X _21025_/X VGND VGND VPWR VPWR _21027_/A
+ sky130_fd_sc_hd__a41o_4
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23008__B _23008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22898__B1 _24422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22977_ _21546_/X _22974_/Y _22423_/X _22976_/X VGND VGND VPWR VPWR _22977_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19763__B1 _19714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12730_ _12730_/A _12730_/B VGND VGND VPWR VPWR _12732_/B sky130_fd_sc_hd__or2_4
X_24716_ _23664_/CLK _24716_/D HRESETn VGND VGND VPWR VPWR _14683_/A sky130_fd_sc_hd__dfrtp_4
X_21928_ _21159_/A _21928_/B VGND VGND VPWR VPWR _21928_/X sky130_fd_sc_hd__or2_4
XANTENNA__16577__B1 _16246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12661_ _12637_/X _12659_/X _12660_/X VGND VGND VPWR VPWR _25068_/D sky130_fd_sc_hd__and3_4
XFILLER_76_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21859_ _22226_/A _21858_/X _16371_/Y _20757_/X VGND VGND VPWR VPWR _21859_/X sky130_fd_sc_hd__o22a_4
XFILLER_128_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24647_ _24644_/CLK _24647_/D HRESETn VGND VGND VPWR VPWR _13717_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_19_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _13663_/A VGND VGND VPWR VPWR _11612_/X sky130_fd_sc_hd__buf_2
X_14400_ _14385_/A _14384_/X VGND VGND VPWR VPWR _14400_/Y sky130_fd_sc_hd__nand2_4
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _24519_/Q VGND VGND VPWR VPWR _12592_/Y sky130_fd_sc_hd__inv_2
X_15380_ _24593_/Q VGND VGND VPWR VPWR _22212_/A sky130_fd_sc_hd__inv_2
XANTENNA__16329__B1 _15484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11989__B _11956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19556__A2_N _19555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24578_ _25183_/CLK _24578_/D HRESETn VGND VGND VPWR VPWR _14432_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ _11539_/Y _11521_/X _11540_/X _11542_/X VGND VGND VPWR VPWR _25217_/D sky130_fd_sc_hd__a2bb2o_4
X_14331_ _14320_/Y VGND VGND VPWR VPWR _14331_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_49_0_HCLK clkbuf_7_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_99_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23529_ _23537_/CLK _18892_/X VGND VGND VPWR VPWR _23529_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21070__A2_N _22322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ _24801_/Q VGND VGND VPWR VPWR _14262_/Y sky130_fd_sc_hd__inv_2
X_17050_ _24058_/Q _17051_/B VGND VGND VPWR VPWR _17050_/X sky130_fd_sc_hd__or2_4
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24287__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13213_ _13309_/A _23378_/Q VGND VGND VPWR VPWR _13213_/X sky130_fd_sc_hd__or2_4
X_16001_ _24360_/Q VGND VGND VPWR VPWR _16001_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15477__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14193_ _20195_/A VGND VGND VPWR VPWR _20193_/A sky130_fd_sc_hd__inv_2
XFILLER_136_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24216__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13144_ _13182_/A _13144_/B VGND VGND VPWR VPWR _13144_/X sky130_fd_sc_hd__or2_4
XFILLER_3_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21085__A2_N _21083_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17692__A _14569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13075_ _13075_/A VGND VGND VPWR VPWR _13203_/A sky130_fd_sc_hd__buf_2
X_17952_ _17821_/A _17952_/B VGND VGND VPWR VPWR _17952_/X sky130_fd_sc_hd__or2_4
XANTENNA__21926__B _21924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12026_ _23795_/Q _12014_/B _12025_/Y VGND VGND VPWR VPWR _12026_/X sky130_fd_sc_hd__o21a_4
X_16903_ _16890_/A _16900_/B _16903_/C VGND VGND VPWR VPWR _16903_/X sky130_fd_sc_hd__and3_4
XFILLER_78_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17883_ _17947_/A _17883_/B _17883_/C VGND VGND VPWR VPWR _17891_/B sky130_fd_sc_hd__or3_4
XANTENNA__15068__B1 _15027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22103__A _20966_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20061__B1 _19424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19622_ _19530_/X _19282_/B _19236_/X VGND VGND VPWR VPWR _19623_/A sky130_fd_sc_hd__or3_4
X_16834_ _16832_/Y _16778_/Y _16834_/C _16834_/D VGND VGND VPWR VPWR _16834_/X sky130_fd_sc_hd__or4_4
XFILLER_76_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14815__B1 _14990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23851__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19553_ _18018_/X _18025_/D _19531_/X VGND VGND VPWR VPWR _19554_/A sky130_fd_sc_hd__or3_4
X_16765_ _16765_/A VGND VGND VPWR VPWR _16765_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22889__B1 _12089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13977_ _24888_/Q _13928_/B _24888_/Q _13928_/B VGND VGND VPWR VPWR _13977_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25075__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18504_ _18504_/A _18504_/B _18503_/X VGND VGND VPWR VPWR _23830_/D sky130_fd_sc_hd__and3_4
XFILLER_46_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16754__A1_N _15892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15716_ _15716_/A VGND VGND VPWR VPWR _15717_/B sky130_fd_sc_hd__inv_2
XANTENNA__15940__A _22783_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12928_ _22769_/A _12931_/B VGND VGND VPWR VPWR _12929_/C sky130_fd_sc_hd__or2_4
X_19484_ _23319_/Q VGND VGND VPWR VPWR _19484_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25004__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16696_ _16689_/X _16691_/X _16694_/X _16696_/D VGND VGND VPWR VPWR _16717_/B sky130_fd_sc_hd__or4_4
X_18435_ _18518_/A _18515_/A _18432_/X _18434_/X VGND VGND VPWR VPWR _18436_/B sky130_fd_sc_hd__or4_4
X_15647_ _15460_/X VGND VGND VPWR VPWR _15647_/X sky130_fd_sc_hd__buf_2
X_12859_ _12858_/X _24432_/Q _25006_/Q _12826_/Y VGND VGND VPWR VPWR _12859_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16139__A1_N _16133_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18366_ _16457_/A _23820_/Q _16457_/Y _18535_/A VGND VGND VPWR VPWR _18366_/X sky130_fd_sc_hd__o22a_4
X_15578_ _15414_/A _15578_/B VGND VGND VPWR VPWR _15578_/X sky130_fd_sc_hd__or2_4
X_17317_ _17262_/Y _17413_/A _17317_/C _17317_/D VGND VGND VPWR VPWR _17324_/A sky130_fd_sc_hd__or4_4
XFILLER_30_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14529_ _21007_/A VGND VGND VPWR VPWR _14529_/X sky130_fd_sc_hd__buf_2
X_18297_ _18218_/B _18292_/B _18294_/B _18228_/X VGND VGND VPWR VPWR _18298_/A sky130_fd_sc_hd__a211o_4
X_17248_ _25211_/Q _17246_/Y _25217_/Q _17353_/A VGND VGND VPWR VPWR _17248_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15387__A _15358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_6_0_HCLK clkbuf_6_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_17179_ _23675_/Q _17179_/B VGND VGND VPWR VPWR _20385_/B sky130_fd_sc_hd__or2_4
X_20190_ _23777_/Q _20234_/B _20178_/A VGND VGND VPWR VPWR _20191_/B sky130_fd_sc_hd__and3_4
XFILLER_115_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23939__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19634__A1_N _21469_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22900_ _22900_/A _22651_/B VGND VGND VPWR VPWR _22900_/X sky130_fd_sc_hd__and2_4
X_23880_ _24984_/CLK _18126_/X HRESETn VGND VGND VPWR VPWR _18124_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14806__B1 _14703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21852__A _21034_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22831_ _22201_/A _22816_/X _22819_/X _22825_/X _22830_/X VGND VGND VPWR VPWR _22831_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22762_ _22597_/A _22761_/X VGND VGND VPWR VPWR _22762_/X sky130_fd_sc_hd__and2_4
XFILLER_25_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21713_ _20837_/X _21707_/X _21708_/X _21175_/X _21712_/Y VGND VGND VPWR VPWR _21713_/X
+ sky130_fd_sc_hd__a32o_4
X_24501_ _23949_/CLK _15646_/X HRESETn VGND VGND VPWR VPWR _20739_/B sky130_fd_sc_hd__dfrtp_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22693_ _24345_/Q _22549_/A _22581_/X VGND VGND VPWR VPWR _22693_/X sky130_fd_sc_hd__o21a_4
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16574__A3 HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24798__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21644_ _21644_/A _21181_/A VGND VGND VPWR VPWR _21644_/X sky130_fd_sc_hd__and2_4
X_24432_ _24432_/CLK _15800_/X HRESETn VGND VGND VPWR VPWR _24432_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24727__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20658__A2 _20552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24363_ _24425_/CLK _15996_/X HRESETn VGND VGND VPWR VPWR _24363_/Q sky130_fd_sc_hd__dfrtp_4
X_21575_ _23731_/Q VGND VGND VPWR VPWR _21575_/Y sky130_fd_sc_hd__inv_2
X_23314_ _23313_/CLK _23314_/D VGND VGND VPWR VPWR _23314_/Q sky130_fd_sc_hd__dfxtp_4
X_20526_ _20511_/X _20525_/Y _24608_/Q _20515_/X VGND VGND VPWR VPWR _20526_/X sky130_fd_sc_hd__a2bb2o_4
X_24294_ _24319_/CLK _16206_/X HRESETn VGND VGND VPWR VPWR _24294_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24380__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23245_ _23278_/CLK _23245_/D VGND VGND VPWR VPWR _23245_/Q sky130_fd_sc_hd__dfxtp_4
X_20457_ _13506_/C VGND VGND VPWR VPWR _20457_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23176_ _25112_/CLK _23176_/D VGND VGND VPWR VPWR _23176_/Q sky130_fd_sc_hd__dfxtp_4
X_20388_ _20388_/A VGND VGND VPWR VPWR _20388_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20931__A _20931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22127_ _22155_/A _22126_/X _21986_/X _24509_/Q _21987_/X VGND VGND VPWR VPWR _22127_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21746__B _15639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22058_ _21675_/A _22056_/X _22057_/X VGND VGND VPWR VPWR _22058_/X sky130_fd_sc_hd__and3_4
XFILLER_43_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13900_ _13908_/A _13900_/B VGND VGND VPWR VPWR _13900_/X sky130_fd_sc_hd__and2_4
X_21009_ _21009_/A _19837_/Y VGND VGND VPWR VPWR _21010_/C sky130_fd_sc_hd__or2_4
X_14880_ _14880_/A _14879_/X VGND VGND VPWR VPWR _14995_/A sky130_fd_sc_hd__or2_4
XANTENNA__22858__A _22858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13831_ _13824_/X _13825_/X _13831_/C _13830_/X VGND VGND VPWR VPWR _13869_/D sky130_fd_sc_hd__or4_4
XFILLER_112_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16856__A _16774_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16550_ _16548_/Y _16542_/X _16211_/X _16549_/X VGND VGND VPWR VPWR _24161_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21481__B _19698_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19232__A _18711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13762_ _13770_/A _13776_/B _13776_/C _13762_/D VGND VGND VPWR VPWR _13763_/A sky130_fd_sc_hd__or4_4
Xclkbuf_5_12_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_15501_ HWDATA[13] VGND VGND VPWR VPWR _15501_/X sky130_fd_sc_hd__buf_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12713_ _12554_/X _12710_/D VGND VGND VPWR VPWR _12714_/B sky130_fd_sc_hd__or2_4
X_16481_ _16493_/A VGND VGND VPWR VPWR _16481_/X sky130_fd_sc_hd__buf_2
X_13693_ _13682_/Y VGND VGND VPWR VPWR _13693_/X sky130_fd_sc_hd__buf_2
X_18220_ _18242_/A _18242_/B _18201_/X _18219_/X VGND VGND VPWR VPWR _18221_/C sky130_fd_sc_hd__or4_4
XANTENNA__13280__A _13092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15432_ _15431_/X VGND VGND VPWR VPWR _15432_/X sky130_fd_sc_hd__buf_2
X_12644_ _12565_/Y _12554_/X _12609_/Y _12644_/D VGND VGND VPWR VPWR _12644_/X sky130_fd_sc_hd__or4_4
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24468__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18151_ _16063_/A _23869_/Q _16063_/Y _18242_/B VGND VGND VPWR VPWR _18151_/X sky130_fd_sc_hd__o22a_4
XFILLER_129_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ _24509_/Q VGND VGND VPWR VPWR _12575_/Y sky130_fd_sc_hd__inv_2
X_15363_ _15363_/A VGND VGND VPWR VPWR _15363_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21846__B2 _20900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17102_ _17097_/A _17097_/B _17083_/X _17099_/B VGND VGND VPWR VPWR _17102_/X sky130_fd_sc_hd__a211o_4
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14314_ _23650_/Q VGND VGND VPWR VPWR _14315_/C sky130_fd_sc_hd__inv_2
X_11526_ _11524_/Y _11521_/X _11525_/X _11521_/X VGND VGND VPWR VPWR _11526_/X sky130_fd_sc_hd__a2bb2o_4
X_18082_ _13011_/X _18081_/X _13011_/X _18081_/X VGND VGND VPWR VPWR _23893_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15294_ _15294_/A VGND VGND VPWR VPWR _15294_/Y sky130_fd_sc_hd__inv_2
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17033_ _16966_/Y _17144_/A VGND VGND VPWR VPWR _17033_/X sky130_fd_sc_hd__or2_4
X_14245_ _14004_/Y _14243_/X _14094_/X _14243_/X VGND VGND VPWR VPWR _14245_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_136_0_HCLK clkbuf_7_68_0_HCLK/X VGND VGND VPWR VPWR _23442_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24050__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14176_ _14165_/B VGND VGND VPWR VPWR _14176_/X sky130_fd_sc_hd__buf_2
XANTENNA__21937__A _21172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_199_0_HCLK clkbuf_7_99_0_HCLK/X VGND VGND VPWR VPWR _24167_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_113_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15289__B1 _14304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13127_ _13127_/A _20140_/A VGND VGND VPWR VPWR _13129_/B sky130_fd_sc_hd__or2_4
X_18984_ _23496_/Q VGND VGND VPWR VPWR _18984_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22023__A1 _22223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13058_ _11733_/A VGND VGND VPWR VPWR _13073_/A sky130_fd_sc_hd__buf_2
X_17935_ _17935_/A _17935_/B VGND VGND VPWR VPWR _17936_/C sky130_fd_sc_hd__or2_4
XFILLER_97_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12009_ _25139_/Q VGND VGND VPWR VPWR _12054_/A sky130_fd_sc_hd__inv_2
XANTENNA__13455__A _13454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17866_ _17898_/A _17866_/B _17865_/X VGND VGND VPWR VPWR _17874_/B sky130_fd_sc_hd__or3_4
XFILLER_94_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12392__A1_N _12391_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16817_ _16817_/A VGND VGND VPWR VPWR _16920_/A sky130_fd_sc_hd__inv_2
X_19605_ _19602_/Y _19596_/X _19603_/X _19604_/X VGND VGND VPWR VPWR _23276_/D sky130_fd_sc_hd__a2bb2o_4
X_17797_ _17796_/X _23524_/Q VGND VGND VPWR VPWR _17798_/C sky130_fd_sc_hd__or2_4
XANTENNA__22487__B _22188_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19536_ _23301_/Q VGND VGND VPWR VPWR _19536_/Y sky130_fd_sc_hd__inv_2
X_16748_ _16747_/Y VGND VGND VPWR VPWR _16748_/X sky130_fd_sc_hd__buf_2
XANTENNA__20337__A1 _20331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19467_ _19467_/A VGND VGND VPWR VPWR _19467_/Y sky130_fd_sc_hd__inv_2
X_16679_ _14564_/X _14598_/Y _16678_/X _14597_/X VGND VGND VPWR VPWR _16679_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24891__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18418_ _18416_/Y _18470_/A VGND VGND VPWR VPWR _18437_/C sky130_fd_sc_hd__or2_4
X_19398_ _19394_/Y _19397_/X _19329_/X _19397_/X VGND VGND VPWR VPWR _19398_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24820__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21837__A1 _20750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18349_ _23823_/Q VGND VGND VPWR VPWR _18425_/A sky130_fd_sc_hd__inv_2
XFILLER_124_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21837__B2 _21836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24138__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21360_ _11941_/X VGND VGND VPWR VPWR _22548_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_32_0_HCLK clkbuf_6_16_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_65_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20311_ _18616_/B _20310_/Y _20315_/C VGND VGND VPWR VPWR _20311_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_95_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_95_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21291_ _21291_/A _20749_/X VGND VGND VPWR VPWR _21296_/B sky130_fd_sc_hd__or2_4
XANTENNA__12534__A _12534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23030_ _22997_/A _23030_/B _23030_/C _23029_/Y VGND VGND VPWR VPWR _23030_/X sky130_fd_sc_hd__or4_4
X_20242_ _20254_/A _20241_/Y VGND VGND VPWR VPWR _20243_/C sky130_fd_sc_hd__and2_4
XFILLER_131_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16646__A1_N _14751_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20173_ _20173_/A _20194_/A _20196_/A _20172_/X VGND VGND VPWR VPWR _20173_/X sky130_fd_sc_hd__or4_4
XANTENNA__21566__B _20818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23773__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_1_0_HCLK clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_24981_ _24984_/CLK _13373_/X HRESETn VGND VGND VPWR VPWR _11890_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19966__B1 _19392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23702__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23932_ _24735_/CLK _17768_/X HRESETn VGND VGND VPWR VPWR _23932_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23863_ _23859_/CLK _23863_/D HRESETn VGND VGND VPWR VPWR _23863_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15580__A _15741_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24979__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22814_ _24492_/Q _20757_/A VGND VGND VPWR VPWR _22814_/X sky130_fd_sc_hd__or2_4
XFILLER_44_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23794_ _23796_/CLK _20694_/X HRESETn VGND VGND VPWR VPWR _23794_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24908__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22745_ _24116_/Q _22745_/B VGND VGND VPWR VPWR _22745_/X sky130_fd_sc_hd__or2_4
XANTENNA__15204__B1 _15147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14196__A _16231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18891__A _18876_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18941__B2 _18935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22676_ _24415_/Q _22281_/X _22558_/X _22675_/X VGND VGND VPWR VPWR _22676_/X sky130_fd_sc_hd__a211o_4
XFILLER_129_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20926__A _20926_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24561__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21627_ _21623_/X _21626_/X _18048_/X VGND VGND VPWR VPWR _21627_/X sky130_fd_sc_hd__o21a_4
X_24415_ _24425_/CLK _24415_/D HRESETn VGND VGND VPWR VPWR _24415_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12360_ _12360_/A VGND VGND VPWR VPWR _12495_/A sky130_fd_sc_hd__buf_2
X_21558_ _17208_/A _21553_/X _21555_/X _21556_/X _21557_/X VGND VGND VPWR VPWR _21558_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24346_ _23872_/CLK _16069_/X HRESETn VGND VGND VPWR VPWR _24346_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20509_ _20513_/B _20502_/X _20508_/X VGND VGND VPWR VPWR _20509_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_5_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12291_ _12265_/C _12298_/A VGND VGND VPWR VPWR _12300_/A sky130_fd_sc_hd__or2_4
X_24277_ _24681_/CLK _16255_/X HRESETn VGND VGND VPWR VPWR _14960_/A sky130_fd_sc_hd__dfrtp_4
X_21489_ _21473_/X _21488_/X _20820_/X VGND VGND VPWR VPWR _21489_/Y sky130_fd_sc_hd__a21oi_4
X_14030_ _20245_/A VGND VGND VPWR VPWR _20239_/A sky130_fd_sc_hd__inv_2
XFILLER_4_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_209_0_HCLK clkbuf_7_104_0_HCLK/X VGND VGND VPWR VPWR _24225_/CLK sky130_fd_sc_hd__clkbuf_1
X_23228_ _23246_/CLK _19744_/X VGND VGND VPWR VPWR _19742_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_107_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18457__B1 _18449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19227__A _11635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23159_ _25106_/CLK _19923_/X VGND VGND VPWR VPWR _23159_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_122_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22005__B2 _21570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15981_ _15981_/A VGND VGND VPWR VPWR _15981_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15691__B1 _22373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17720_ _17729_/A VGND VGND VPWR VPWR _17721_/A sky130_fd_sc_hd__buf_2
XANTENNA__24803__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14932_ _14893_/X _14932_/B _14918_/X _14931_/X VGND VGND VPWR VPWR _14974_/A sky130_fd_sc_hd__or4_4
XANTENNA__24866__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17651_ _17651_/A VGND VGND VPWR VPWR _21335_/A sky130_fd_sc_hd__buf_2
X_14863_ _14841_/X _14848_/X _14855_/X _14862_/X VGND VGND VPWR VPWR _14863_/X sky130_fd_sc_hd__or4_4
XFILLER_91_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16602_ _16584_/A VGND VGND VPWR VPWR _16602_/X sky130_fd_sc_hd__buf_2
XFILLER_90_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13814_ _13869_/A VGND VGND VPWR VPWR _13852_/A sky130_fd_sc_hd__buf_2
XFILLER_21_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17582_ _17547_/X _17580_/X _17581_/X VGND VGND VPWR VPWR _23955_/D sky130_fd_sc_hd__and3_4
X_14794_ _14794_/A _14794_/B _14784_/X _14794_/D VGND VGND VPWR VPWR _14794_/X sky130_fd_sc_hd__or4_4
XFILLER_91_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19321_ _13277_/B VGND VGND VPWR VPWR _19321_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24649__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16533_ _16532_/Y _16530_/X _16451_/X _16530_/X VGND VGND VPWR VPWR _16533_/X sky130_fd_sc_hd__a2bb2o_4
X_13745_ _13745_/A _13745_/B _13737_/Y _13745_/D VGND VGND VPWR VPWR _13792_/B sky130_fd_sc_hd__and4_4
XFILLER_71_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19252_ _19250_/Y _19251_/X _11857_/X _19251_/X VGND VGND VPWR VPWR _19252_/X sky130_fd_sc_hd__a2bb2o_4
X_16464_ _24194_/Q VGND VGND VPWR VPWR _16464_/Y sky130_fd_sc_hd__inv_2
X_13676_ _23688_/Q VGND VGND VPWR VPWR _13677_/C sky130_fd_sc_hd__inv_2
XANTENNA__20836__A _20820_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18203_ _23860_/Q VGND VGND VPWR VPWR _18203_/Y sky130_fd_sc_hd__inv_2
X_15415_ _16475_/B VGND VGND VPWR VPWR _15415_/Y sky130_fd_sc_hd__inv_2
X_12627_ _25065_/Q _12615_/Y _12737_/A _15630_/A VGND VGND VPWR VPWR _12627_/X sky130_fd_sc_hd__a2bb2o_4
X_19183_ _19181_/Y _19182_/X _19115_/X _19182_/X VGND VGND VPWR VPWR _23425_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16395_ _16401_/A VGND VGND VPWR VPWR _16395_/X sky130_fd_sc_hd__buf_2
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24231__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18134_ _23851_/Q VGND VGND VPWR VPWR _18318_/A sky130_fd_sc_hd__inv_2
X_15346_ _22753_/A _15340_/X _11555_/X _15345_/X VGND VGND VPWR VPWR _24607_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21295__A2 _21292_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12558_ _12648_/A _12556_/Y _12679_/C _24528_/Q VGND VGND VPWR VPWR _12558_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_19_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11509_ _24622_/Q VGND VGND VPWR VPWR _15314_/A sky130_fd_sc_hd__inv_2
X_18065_ _11755_/A _18065_/B _18065_/C _18064_/X VGND VGND VPWR VPWR _19801_/B sky130_fd_sc_hd__and4_4
XFILLER_8_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15277_ _15275_/Y _15272_/X _14236_/X _15276_/X VGND VGND VPWR VPWR _15277_/X sky130_fd_sc_hd__a2bb2o_4
X_12489_ _12489_/A _12489_/B VGND VGND VPWR VPWR _12490_/C sky130_fd_sc_hd__or2_4
X_17016_ _16202_/Y _16961_/A _16210_/Y _24030_/Q VGND VGND VPWR VPWR _17016_/X sky130_fd_sc_hd__a2bb2o_4
X_14228_ _16369_/A VGND VGND VPWR VPWR _14228_/X sky130_fd_sc_hd__buf_2
XANTENNA__22244__A1 _22501_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12159__A2_N _12075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14159_ _18111_/C VGND VGND VPWR VPWR _14159_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18967_ _11755_/A _23894_/Q _11729_/X VGND VGND VPWR VPWR _20134_/C sky130_fd_sc_hd__or3_4
XANTENNA__25090__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13185__A _11751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15682__B1 _11570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17918_ _17918_/A _17918_/B _17918_/C VGND VGND VPWR VPWR _17922_/B sky130_fd_sc_hd__and3_4
XFILLER_100_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18898_ _19946_/C _19167_/B _18920_/A _19189_/B VGND VGND VPWR VPWR _18898_/X sky130_fd_sc_hd__or4_4
XFILLER_66_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22498__A _15363_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17849_ _17881_/A _23146_/Q VGND VGND VPWR VPWR _17850_/C sky130_fd_sc_hd__or2_4
XFILLER_6_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20860_ _16125_/Y _21093_/B _21882_/A _20859_/X VGND VGND VPWR VPWR _20863_/B sky130_fd_sc_hd__a211o_4
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19519_ _21676_/B _19516_/X _19452_/X _19516_/X VGND VGND VPWR VPWR _23307_/D sky130_fd_sc_hd__a2bb2o_4
X_20791_ _21448_/B _20790_/X _24392_/Q _11940_/Y VGND VGND VPWR VPWR _20791_/X sky130_fd_sc_hd__o22a_4
XFILLER_35_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24319__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22530_ _22610_/A VGND VGND VPWR VPWR _22530_/X sky130_fd_sc_hd__buf_2
XANTENNA__15737__A1 _15582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20746__A _20745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22461_ _20909_/X _22458_/X _22459_/X _11579_/A _22460_/X VGND VGND VPWR VPWR _22461_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_22_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14744__A _14744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21412_ _22444_/B _21411_/X _21046_/X _25193_/Q _21047_/X VGND VGND VPWR VPWR _21413_/A
+ sky130_fd_sc_hd__a32o_4
X_24200_ _24197_/CLK _24200_/D HRESETn VGND VGND VPWR VPWR _16448_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25180_ _24847_/CLK _11816_/Y HRESETn VGND VGND VPWR VPWR _25180_/Q sky130_fd_sc_hd__dfrtp_4
X_22392_ _13360_/A _22391_/X _22251_/X _24558_/Q _21059_/X VGND VGND VPWR VPWR _22392_/X
+ sky130_fd_sc_hd__a32o_4
X_24131_ _24101_/CLK _16611_/X HRESETn VGND VGND VPWR VPWR _14836_/A sky130_fd_sc_hd__dfrtp_4
X_21343_ _21155_/A _21343_/B _21342_/X VGND VGND VPWR VPWR _21343_/X sky130_fd_sc_hd__and3_4
XANTENNA__23954__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24062_ _24618_/CLK _24062_/D HRESETn VGND VGND VPWR VPWR _24062_/Q sky130_fd_sc_hd__dfrtp_4
X_21274_ _24192_/Q _22444_/B VGND VGND VPWR VPWR _21274_/X sky130_fd_sc_hd__or2_4
XFILLER_116_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25178__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23013_ _23013_/A _22245_/A VGND VGND VPWR VPWR _23013_/X sky130_fd_sc_hd__and2_4
X_20225_ _23772_/Q _20225_/B VGND VGND VPWR VPWR _20225_/X sky130_fd_sc_hd__and2_4
XANTENNA__22786__A2 _22259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25107__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_182_0_HCLK clkbuf_7_91_0_HCLK/X VGND VGND VPWR VPWR _24483_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20156_ _14206_/A _20193_/C VGND VGND VPWR VPWR _20156_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_39_0_HCLK clkbuf_8_39_0_HCLK/A VGND VGND VPWR VPWR _25002_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22538__A2 _22536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17790__A _17918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20087_ _20086_/Y _20082_/X _19610_/A _20082_/X VGND VGND VPWR VPWR _20087_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20549__A1 _20413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24964_ _24013_/CLK _13547_/X HRESETn VGND VGND VPWR VPWR _24964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20549__B2 _20465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12430__C _12401_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23915_ _24928_/CLK _17997_/X HRESETn VGND VGND VPWR VPWR _23915_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22201__A _22201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24895_ _24884_/CLK _24895_/D HRESETn VGND VGND VPWR VPWR _24895_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11860_ _19617_/A VGND VGND VPWR VPWR _11860_/X sky130_fd_sc_hd__buf_2
XANTENNA__23016__B _22857_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23846_ _23845_/CLK _18335_/X HRESETn VGND VGND VPWR VPWR _18334_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24742__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11791_ _11771_/Y VGND VGND VPWR VPWR _11809_/B sky130_fd_sc_hd__buf_2
X_20989_ _21012_/A _19505_/Y VGND VGND VPWR VPWR _20991_/B sky130_fd_sc_hd__or2_4
X_23777_ _23668_/CLK _20194_/X HRESETn VGND VGND VPWR VPWR _23777_/Q sky130_fd_sc_hd__dfrtp_4
X_13530_ _23731_/Q _13529_/X VGND VGND VPWR VPWR _13531_/B sky130_fd_sc_hd__or2_4
X_22728_ _16330_/Y _21896_/X _16068_/Y _22549_/X VGND VGND VPWR VPWR _22728_/X sky130_fd_sc_hd__o22a_4
X_13461_ _11507_/X _13460_/X _13461_/C _11726_/Y VGND VGND VPWR VPWR _13461_/X sky130_fd_sc_hd__or4_4
X_22659_ _22651_/X _22659_/B _22655_/X _22658_/X VGND VGND VPWR VPWR _22659_/X sky130_fd_sc_hd__or4_4
X_15200_ _15108_/C _15216_/A VGND VGND VPWR VPWR _15213_/B sky130_fd_sc_hd__or2_4
X_12412_ _12412_/A _12412_/B _12412_/C _12412_/D VGND VGND VPWR VPWR _12413_/D sky130_fd_sc_hd__or4_4
X_16180_ _16176_/Y _16178_/X _16179_/X _16178_/X VGND VGND VPWR VPWR _24305_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21277__A2 _22154_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13392_ _24978_/Q _13390_/Y _13391_/X _13388_/B VGND VGND VPWR VPWR _13392_/X sky130_fd_sc_hd__a211o_4
XFILLER_16_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15131_ _24679_/Q _15130_/Y VGND VGND VPWR VPWR _15131_/X sky130_fd_sc_hd__or2_4
X_12343_ _12432_/A _24496_/Q _12433_/A _12342_/Y VGND VGND VPWR VPWR _12351_/B sky130_fd_sc_hd__o22a_4
XANTENNA__17965__A _17716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24329_ _23852_/CLK _24329_/D HRESETn VGND VGND VPWR VPWR _24329_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23695__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12274_ _12178_/C _12276_/B _12273_/Y VGND VGND VPWR VPWR _12274_/X sky130_fd_sc_hd__o21a_4
X_15062_ _15064_/B VGND VGND VPWR VPWR _15063_/B sky130_fd_sc_hd__inv_2
XANTENNA__17684__B _17684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14013_ _14013_/A _14013_/B VGND VGND VPWR VPWR _15407_/A sky130_fd_sc_hd__or2_4
XANTENNA__23624__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19870_ _21780_/B _19864_/X _19821_/X _19869_/X VGND VGND VPWR VPWR _23180_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18821_ _13226_/B VGND VGND VPWR VPWR _18821_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18850__B1 _18662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18752_ _18752_/A VGND VGND VPWR VPWR _18752_/X sky130_fd_sc_hd__buf_2
XFILLER_136_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15964_ _15963_/Y _15961_/X _11581_/X _15961_/X VGND VGND VPWR VPWR _15964_/X sky130_fd_sc_hd__a2bb2o_4
X_17703_ _17699_/X _17702_/X _14564_/X VGND VGND VPWR VPWR _17703_/X sky130_fd_sc_hd__o21a_4
X_14915_ _14915_/A VGND VGND VPWR VPWR _15108_/C sky130_fd_sc_hd__inv_2
X_18683_ _18681_/Y _18682_/X _16671_/X _18682_/X VGND VGND VPWR VPWR _18683_/X sky130_fd_sc_hd__a2bb2o_4
X_15895_ _15892_/Y _15893_/X _15894_/X _15893_/X VGND VGND VPWR VPWR _15895_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22111__A _20975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17634_ _17634_/A VGND VGND VPWR VPWR _17634_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17205__A _16376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14846_ _14757_/Y VGND VGND VPWR VPWR _15019_/B sky130_fd_sc_hd__buf_2
XFILLER_90_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24483__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17565_ _17565_/A VGND VGND VPWR VPWR _17565_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14777_ _14777_/A VGND VGND VPWR VPWR _14777_/Y sky130_fd_sc_hd__inv_2
X_11989_ _15271_/A _11956_/X VGND VGND VPWR VPWR _11990_/A sky130_fd_sc_hd__nor2_4
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22162__B1 _20744_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12349__A _12349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19304_ _19304_/A VGND VGND VPWR VPWR _19304_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24412__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16516_ _16515_/Y _16511_/X _16179_/X _16511_/X VGND VGND VPWR VPWR _24174_/D sky130_fd_sc_hd__a2bb2o_4
X_13728_ _13728_/A VGND VGND VPWR VPWR _13728_/X sky130_fd_sc_hd__buf_2
X_17496_ _22434_/A VGND VGND VPWR VPWR _17497_/B sky130_fd_sc_hd__inv_2
XANTENNA__20016__A2_N _20015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19235_ _18031_/B VGND VGND VPWR VPWR _19282_/B sky130_fd_sc_hd__buf_2
X_16447_ _16445_/Y _16446_/X _16100_/X _16446_/X VGND VGND VPWR VPWR _24201_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13659_ _22271_/A _13657_/X _13658_/X _13657_/X VGND VGND VPWR VPWR _24935_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19166_ _23430_/Q VGND VGND VPWR VPWR _19166_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18669__B1 _17199_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16378_ _16378_/A VGND VGND VPWR VPWR _16378_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18117_ _23883_/Q VGND VGND VPWR VPWR _18117_/Y sky130_fd_sc_hd__inv_2
X_15329_ _15329_/A VGND VGND VPWR VPWR _15329_/Y sky130_fd_sc_hd__inv_2
X_19097_ _23455_/Q VGND VGND VPWR VPWR _19097_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23009__A3 _22839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18048_ _18047_/Y VGND VGND VPWR VPWR _18048_/X sky130_fd_sc_hd__buf_2
XANTENNA__15498__A3 _15497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13908__A _13908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25200__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20010_ _20010_/A VGND VGND VPWR VPWR _20010_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_255_0_HCLK clkbuf_8_255_0_HCLK/A VGND VGND VPWR VPWR _24671_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21440__A2 _13357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19999_ _19998_/Y _19996_/X _15520_/X _19996_/X VGND VGND VPWR VPWR _23131_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23762__D _23762_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22659__C _22655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21961_ _21229_/A _19578_/Y VGND VGND VPWR VPWR _21961_/X sky130_fd_sc_hd__or2_4
XANTENNA__14739__A _24711_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22940__A2 _22536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23700_ _24162_/CLK _20441_/Y HRESETn VGND VGND VPWR VPWR _20438_/A sky130_fd_sc_hd__dfrtp_4
X_20912_ _22014_/B VGND VGND VPWR VPWR _21860_/B sky130_fd_sc_hd__buf_2
X_21892_ _14230_/Y _20818_/X _24806_/Q _21868_/B VGND VGND VPWR VPWR _21892_/X sky130_fd_sc_hd__a2bb2o_4
X_24680_ _24681_/CLK _24680_/D HRESETn VGND VGND VPWR VPWR _24680_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11692__B2 _11691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21860__A _14887_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _11725_/X VGND VGND VPWR VPWR _20844_/B sky130_fd_sc_hd__buf_2
XPHY_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23631_ _23641_/CLK _23631_/D HRESETn VGND VGND VPWR VPWR _23631_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24153__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20774_ _21990_/A VGND VGND VPWR VPWR _21850_/A sky130_fd_sc_hd__buf_2
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23562_ _23563_/CLK _18796_/X VGND VGND VPWR VPWR _17861_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22513_ _22832_/C VGND VGND VPWR VPWR _22661_/C sky130_fd_sc_hd__buf_2
XFILLER_52_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23493_ _23493_/CLK _18994_/X VGND VGND VPWR VPWR _23493_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22444_ _24107_/Q _22444_/B VGND VGND VPWR VPWR _22444_/X sky130_fd_sc_hd__or2_4
X_22375_ _20747_/X _22372_/Y _20815_/X _22374_/X VGND VGND VPWR VPWR _22375_/X sky130_fd_sc_hd__a2bb2o_4
X_25163_ _24623_/CLK _25163_/D HRESETn VGND VGND VPWR VPWR _25163_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_129_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21326_ _21352_/A _21326_/B VGND VGND VPWR VPWR _21326_/X sky130_fd_sc_hd__or2_4
XANTENNA__12604__A2_N _24515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24114_ _24112_/CLK _24114_/D HRESETn VGND VGND VPWR VPWR _24114_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22208__B2 _22931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25094_ _25097_/CLK _12455_/Y HRESETn VGND VGND VPWR VPWR _25094_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21100__A _14754_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21257_ _21257_/A _20780_/A VGND VGND VPWR VPWR _21257_/X sky130_fd_sc_hd__and2_4
XFILLER_11_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19085__B1 _19041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24045_ _24308_/CLK _24045_/D HRESETn VGND VGND VPWR VPWR _24045_/Q sky130_fd_sc_hd__dfrtp_4
X_20208_ _20207_/X VGND VGND VPWR VPWR _20208_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21188_ _21188_/A _21187_/X VGND VGND VPWR VPWR _21188_/X sky130_fd_sc_hd__and2_4
XFILLER_77_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24994__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20139_ _20138_/Y _20136_/X _19421_/X _20136_/X VGND VGND VPWR VPWR _20139_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21982__A3 _21981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24923__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12961_ _12961_/A VGND VGND VPWR VPWR _25019_/D sky130_fd_sc_hd__inv_2
X_24947_ _24957_/CLK _24947_/D HRESETn VGND VGND VPWR VPWR _11683_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_46_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22392__B1 _24558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14700_ _14997_/A VGND VGND VPWR VPWR _14881_/A sky130_fd_sc_hd__inv_2
X_11912_ _11910_/A _11909_/X _11910_/Y _11911_/Y VGND VGND VPWR VPWR _11916_/C sky130_fd_sc_hd__o22a_4
XFILLER_46_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15680_ _15666_/A VGND VGND VPWR VPWR _15680_/X sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_5_15_0_HCLK_A clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12892_ _12915_/C _12867_/X VGND VGND VPWR VPWR _12892_/X sky130_fd_sc_hd__and2_4
X_24878_ _23676_/CLK _14031_/X HRESETn VGND VGND VPWR VPWR _20245_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_22_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14631_ _14617_/C _14631_/B VGND VGND VPWR VPWR _14631_/Y sky130_fd_sc_hd__nor2_4
X_11843_ _19607_/A VGND VGND VPWR VPWR _11843_/Y sky130_fd_sc_hd__inv_2
X_23829_ _23830_/CLK _23829_/D HRESETn VGND VGND VPWR VPWR _23829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17350_ _17306_/Y _17255_/Y _17305_/Y _17358_/B VGND VGND VPWR VPWR _17353_/B sky130_fd_sc_hd__or4_4
X_14562_ _17739_/A _14561_/X _17739_/A _14561_/X VGND VGND VPWR VPWR _14562_/X sky130_fd_sc_hd__a2bb2o_4
X_11774_ _11795_/B VGND VGND VPWR VPWR _11774_/Y sky130_fd_sc_hd__inv_2
X_16301_ _16301_/A _22230_/A VGND VGND VPWR VPWR _16306_/B sky130_fd_sc_hd__or2_4
X_13513_ _20534_/A _13512_/X VGND VGND VPWR VPWR _13513_/X sky130_fd_sc_hd__or2_4
XFILLER_109_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17281_ _11579_/Y _17310_/A _11579_/Y _17310_/A VGND VGND VPWR VPWR _17282_/D sky130_fd_sc_hd__a2bb2o_4
X_14493_ _14493_/A VGND VGND VPWR VPWR _14493_/X sky130_fd_sc_hd__buf_2
XFILLER_105_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19020_ _23483_/Q VGND VGND VPWR VPWR _21663_/B sky130_fd_sc_hd__inv_2
X_16232_ _16235_/B VGND VGND VPWR VPWR _16625_/A sky130_fd_sc_hd__inv_2
X_13444_ _24940_/Q VGND VGND VPWR VPWR _22483_/A sky130_fd_sc_hd__inv_2
XANTENNA__23876__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22447__B2 _22170_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20458__B1 _13506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16163_ _16162_/Y _16158_/X _15765_/X _16158_/X VGND VGND VPWR VPWR _24311_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23805__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13375_ _13374_/Y _13372_/X _11631_/X _13372_/X VGND VGND VPWR VPWR _24980_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25029__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15114_ _15191_/A _14939_/Y _15187_/B VGND VGND VPWR VPWR _15159_/B sky130_fd_sc_hd__or3_4
X_12326_ _22591_/A VGND VGND VPWR VPWR _12326_/Y sky130_fd_sc_hd__inv_2
X_16094_ _22401_/A _16090_/X _16093_/X _16090_/X VGND VGND VPWR VPWR _24337_/D sky130_fd_sc_hd__a2bb2o_4
X_15045_ _15045_/A _15043_/A VGND VGND VPWR VPWR _15046_/C sky130_fd_sc_hd__or2_4
X_19922_ _23159_/Q VGND VGND VPWR VPWR _19922_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19076__B1 _18964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12257_ _12127_/Y _12257_/B VGND VGND VPWR VPWR _12257_/X sky130_fd_sc_hd__or2_4
XFILLER_68_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12188_ _25133_/Q _12188_/B VGND VGND VPWR VPWR _12190_/B sky130_fd_sc_hd__or2_4
X_19853_ _19853_/A VGND VGND VPWR VPWR _19853_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18804_ _17957_/B VGND VGND VPWR VPWR _18804_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_22_0_HCLK clkbuf_8_23_0_HCLK/A VGND VGND VPWR VPWR _24957_/CLK sky130_fd_sc_hd__clkbuf_1
X_16996_ _21124_/A _17160_/A _24294_/Q _17134_/A VGND VGND VPWR VPWR _16996_/X sky130_fd_sc_hd__a2bb2o_4
X_19784_ _19783_/Y _19781_/X _19445_/X _19781_/X VGND VGND VPWR VPWR _19784_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24664__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_85_0_HCLK clkbuf_8_85_0_HCLK/A VGND VGND VPWR VPWR _24904_/CLK sky130_fd_sc_hd__clkbuf_1
X_15947_ _22706_/A VGND VGND VPWR VPWR _15947_/Y sky130_fd_sc_hd__inv_2
X_18735_ _18734_/X VGND VGND VPWR VPWR _18752_/A sky130_fd_sc_hd__inv_2
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22383__B1 _11587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13463__A _13463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18666_ _18968_/A _11761_/A _18666_/C VGND VGND VPWR VPWR _18666_/X sky130_fd_sc_hd__or3_4
X_15878_ _15877_/Y _15873_/X _11594_/X _15873_/X VGND VGND VPWR VPWR _24407_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20933__A1 _15426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16062__B1 _11548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14829_ _14822_/X _14829_/B _14829_/C _14828_/X VGND VGND VPWR VPWR _14829_/X sky130_fd_sc_hd__or4_4
X_17617_ _17487_/Y _17615_/X _17616_/Y VGND VGND VPWR VPWR _23945_/D sky130_fd_sc_hd__o21a_4
X_18597_ _18593_/X _18597_/B _18595_/X _18596_/X VGND VGND VPWR VPWR _18603_/C sky130_fd_sc_hd__or4_4
XANTENNA__16774__A _16774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17548_ _17581_/A _17494_/Y _17586_/A _17492_/X VGND VGND VPWR VPWR _17548_/X sky130_fd_sc_hd__or4_4
X_17479_ _16710_/Y _16733_/Y VGND VGND VPWR VPWR _17505_/B sky130_fd_sc_hd__or2_4
X_19218_ _19212_/Y VGND VGND VPWR VPWR _19218_/X sky130_fd_sc_hd__buf_2
X_20490_ _20499_/C VGND VGND VPWR VPWR _20495_/A sky130_fd_sc_hd__inv_2
X_19149_ _18739_/X VGND VGND VPWR VPWR _19149_/X sky130_fd_sc_hd__buf_2
XANTENNA__22989__A2 _15919_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21839__B _11516_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14708__A2_N _22502_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22160_ _22160_/A _22952_/B VGND VGND VPWR VPWR _22160_/X sky130_fd_sc_hd__or2_4
XANTENNA__22661__D _22660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21111_ _16553_/Y _11529_/A VGND VGND VPWR VPWR _21111_/X sky130_fd_sc_hd__and2_4
XFILLER_12_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15876__B1 _11590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13638__A _15801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22091_ _22084_/A _22091_/B VGND VGND VPWR VPWR _22091_/X sky130_fd_sc_hd__or2_4
XANTENNA__19067__B1 _18953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21042_ _21042_/A VGND VGND VPWR VPWR _21042_/X sky130_fd_sc_hd__buf_2
XFILLER_99_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17617__A1 _17487_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21855__A _21256_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15853__A _24416_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14265__A1_N _14264_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24801_ _24811_/CLK _24801_/D HRESETn VGND VGND VPWR VPWR _24801_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22993_ _15324_/Y _22870_/B VGND VGND VPWR VPWR _22993_/X sky130_fd_sc_hd__and2_4
XFILLER_28_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22374__B1 _24557_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24334__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14851__B2 _14850_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24732_ _23419_/CLK _14603_/X HRESETn VGND VGND VPWR VPWR _24732_/Q sky130_fd_sc_hd__dfrtp_4
X_21944_ _21372_/A _21944_/B _21943_/X VGND VGND VPWR VPWR _21944_/X sky130_fd_sc_hd__and3_4
XANTENNA__12862__B1 _12972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20924__A1 _21553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16053__B1 _15753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20924__B2 _13618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24663_ _24662_/CLK _15192_/X HRESETn VGND VGND VPWR VPWR _15190_/A sky130_fd_sc_hd__dfrtp_4
X_21875_ _24931_/Q _20885_/X VGND VGND VPWR VPWR _21875_/X sky130_fd_sc_hd__or2_4
XPHY_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15800__B1 _24432_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _23493_/CLK _23614_/D VGND VGND VPWR VPWR _23614_/Q sky130_fd_sc_hd__dfxtp_4
X_20826_ _20826_/A VGND VGND VPWR VPWR _20826_/X sky130_fd_sc_hd__buf_2
XPHY_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17499__B _17558_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24594_ _24171_/CLK _15379_/X HRESETn VGND VGND VPWR VPWR _24594_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23545_ _23479_/CLK _23545_/D VGND VGND VPWR VPWR _23545_/Q sky130_fd_sc_hd__dfxtp_4
X_20757_ _20757_/A VGND VGND VPWR VPWR _20757_/X sky130_fd_sc_hd__buf_2
XFILLER_23_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11621__A _11599_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20688_ _20688_/A _20688_/B VGND VGND VPWR VPWR _23785_/D sky130_fd_sc_hd__and2_4
XFILLER_17_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23476_ _23471_/CLK _19043_/X VGND VGND VPWR VPWR _13140_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_137_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25193__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25215_ _24385_/CLK _11549_/X HRESETn VGND VGND VPWR VPWR _11547_/A sky130_fd_sc_hd__dfrtp_4
X_22427_ _22423_/X _22424_/X _22426_/X VGND VGND VPWR VPWR _22457_/B sky130_fd_sc_hd__and3_4
XFILLER_136_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25122__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13160_ _13076_/A VGND VGND VPWR VPWR _13261_/A sky130_fd_sc_hd__buf_2
X_25146_ _24984_/CLK _11993_/X HRESETn VGND VGND VPWR VPWR _11992_/A sky130_fd_sc_hd__dfrtp_4
X_22358_ _22357_/X VGND VGND VPWR VPWR _22358_/Y sky130_fd_sc_hd__inv_2
X_12111_ _24554_/Q VGND VGND VPWR VPWR _12111_/Y sky130_fd_sc_hd__inv_2
X_13091_ _11741_/X VGND VGND VPWR VPWR _13092_/A sky130_fd_sc_hd__buf_2
X_21309_ _24774_/Q _21097_/B VGND VGND VPWR VPWR _21309_/X sky130_fd_sc_hd__and2_4
X_22289_ _16448_/Y _22230_/A _14709_/Y _22547_/A VGND VGND VPWR VPWR _22289_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12452__A _12434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25077_ _25097_/CLK _12521_/X HRESETn VGND VGND VPWR VPWR _25077_/Q sky130_fd_sc_hd__dfrtp_4
X_12042_ _12040_/A _12041_/A _12040_/Y _12041_/Y VGND VGND VPWR VPWR _12045_/C sky130_fd_sc_hd__o22a_4
XANTENNA__21404__A2 _21401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24028_ _24289_/CLK _24028_/D HRESETn VGND VGND VPWR VPWR _21066_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16850_ _16816_/Y _16843_/X _16844_/Y _16849_/X VGND VGND VPWR VPWR _16850_/X sky130_fd_sc_hd__a211o_4
X_15801_ _15801_/A VGND VGND VPWR VPWR _15801_/X sky130_fd_sc_hd__buf_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16292__B1 _16291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16781_ _15862_/A _16780_/A _15862_/Y _16780_/Y VGND VGND VPWR VPWR _16781_/X sky130_fd_sc_hd__o22a_4
X_13993_ _13950_/A _13926_/B _13925_/D _13992_/X VGND VGND VPWR VPWR _13993_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_24_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24075__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18520_ _18515_/A _18515_/B _18475_/X _18517_/B VGND VGND VPWR VPWR _18520_/X sky130_fd_sc_hd__a211o_4
XANTENNA__14842__B2 _24148_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15732_ _24465_/Q _15726_/Y _15722_/C _15731_/X VGND VGND VPWR VPWR _15732_/X sky130_fd_sc_hd__o22a_4
X_12944_ _12809_/Y _12943_/X _12896_/X VGND VGND VPWR VPWR _12944_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__19230__B1 _19207_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20915__A1 _21860_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20678__A1_N _20556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11656__B2 _23914_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20915__B2 _22154_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24004__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18451_ _18451_/A VGND VGND VPWR VPWR _18451_/Y sky130_fd_sc_hd__inv_2
X_15663_ _15658_/X _15647_/X _15468_/X _22975_/A _15661_/X VGND VGND VPWR VPWR _24497_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_2_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12875_ _22258_/A VGND VGND VPWR VPWR _12876_/A sky130_fd_sc_hd__inv_2
XFILLER_73_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17402_ _17315_/A _17401_/Y VGND VGND VPWR VPWR _17402_/X sky130_fd_sc_hd__or2_4
X_14614_ _24727_/Q _14614_/B _14614_/C VGND VGND VPWR VPWR _14615_/A sky130_fd_sc_hd__or3_4
XFILLER_60_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11826_ _11826_/A VGND VGND VPWR VPWR _19597_/A sky130_fd_sc_hd__buf_2
X_18382_ _23818_/Q VGND VGND VPWR VPWR _18421_/B sky130_fd_sc_hd__inv_2
XANTENNA__22668__A1 _21529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15594_ _12560_/Y _15590_/X _11540_/X _15593_/X VGND VGND VPWR VPWR _15594_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22668__B2 _22667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _17237_/Y _17331_/A VGND VGND VPWR VPWR _17334_/C sky130_fd_sc_hd__or2_4
XPHY_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14540_/X _14541_/X _19813_/A VGND VGND VPWR VPWR _14545_/Y sky130_fd_sc_hd__o21ai_4
XPHY_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _11757_/A _23894_/Q VGND VGND VPWR VPWR _17227_/B sky130_fd_sc_hd__and2_4
XPHY_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17544__B1 _17502_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15003__A _15003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17264_ _17264_/A VGND VGND VPWR VPWR _17264_/Y sky130_fd_sc_hd__inv_2
X_14476_ _14429_/X VGND VGND VPWR VPWR _14476_/Y sky130_fd_sc_hd__inv_2
XPHY_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11688_ _23912_/Q VGND VGND VPWR VPWR _11688_/Y sky130_fd_sc_hd__inv_2
X_19003_ _18990_/Y VGND VGND VPWR VPWR _19003_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16215_ _21124_/A VGND VGND VPWR VPWR _16215_/Y sky130_fd_sc_hd__inv_2
X_13427_ _13420_/X _13422_/X _13427_/C _13427_/D VGND VGND VPWR VPWR _13427_/X sky130_fd_sc_hd__or4_4
X_17195_ _23766_/Q _13794_/Y _20733_/A _13794_/A VGND VGND VPWR VPWR _17195_/X sky130_fd_sc_hd__o22a_4
XFILLER_31_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16146_ _16143_/Y _16138_/X _15753_/X _16145_/X VGND VGND VPWR VPWR _16146_/X sky130_fd_sc_hd__a2bb2o_4
X_13358_ _13357_/X VGND VGND VPWR VPWR _13358_/X sky130_fd_sc_hd__buf_2
XANTENNA__19739__A2_N _19738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15858__B1 _15770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12309_ _25076_/Q _12307_/Y _12417_/A _24494_/Q VGND VGND VPWR VPWR _12312_/C sky130_fd_sc_hd__a2bb2o_4
X_16077_ _16075_/Y _16071_/X _15772_/X _16076_/X VGND VGND VPWR VPWR _16077_/X sky130_fd_sc_hd__a2bb2o_4
X_13289_ _13057_/A _13288_/X _24997_/Q _13054_/X VGND VGND VPWR VPWR _24997_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12362__A _12362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24845__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15028_ _15022_/A _15021_/X _15027_/X _15023_/Y VGND VGND VPWR VPWR _15029_/A sky130_fd_sc_hd__a211o_4
X_19905_ _19904_/X VGND VGND VPWR VPWR _19918_/A sky130_fd_sc_hd__inv_2
XANTENNA__21883__A2_N _21882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12068__A1_N SSn_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19836_ _19834_/Y _19831_/X _19835_/X _19831_/X VGND VGND VPWR VPWR _19836_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16283__B1 _15982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19767_ _19767_/A VGND VGND VPWR VPWR _21609_/B sky130_fd_sc_hd__inv_2
X_16979_ _24034_/Q VGND VGND VPWR VPWR _17144_/A sky130_fd_sc_hd__inv_2
X_18718_ _17782_/B VGND VGND VPWR VPWR _18718_/Y sky130_fd_sc_hd__inv_2
X_19698_ _19698_/A VGND VGND VPWR VPWR _19698_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20906__B2 _12063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18649_ _18649_/A VGND VGND VPWR VPWR _18649_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23798__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21660_ _21202_/A _21660_/B _21659_/X VGND VGND VPWR VPWR _21660_/X sky130_fd_sc_hd__and3_4
X_20611_ _20611_/A _20606_/X VGND VGND VPWR VPWR _20611_/X sky130_fd_sc_hd__or2_4
XFILLER_127_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23727__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21591_ _16116_/Y _21591_/B VGND VGND VPWR VPWR _21591_/X sky130_fd_sc_hd__or2_4
XFILLER_71_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12072__B2 _24556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22953__B _22953_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20542_ _20542_/A _20542_/B _13514_/X VGND VGND VPWR VPWR _20542_/X sky130_fd_sc_hd__or3_4
X_23330_ _23313_/CLK _23330_/D VGND VGND VPWR VPWR _23330_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_137_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20473_ _20469_/X VGND VGND VPWR VPWR _20473_/Y sky130_fd_sc_hd__inv_2
X_23261_ _23278_/CLK _19650_/X VGND VGND VPWR VPWR _23261_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25000_ _24998_/CLK _25000_/D HRESETn VGND VGND VPWR VPWR _25000_/Q sky130_fd_sc_hd__dfrtp_4
X_22212_ _22212_/A _22497_/B VGND VGND VPWR VPWR _22212_/X sky130_fd_sc_hd__and2_4
XFILLER_134_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22831__A1 _22201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23192_ _25112_/CLK _19836_/X VGND VGND VPWR VPWR _23192_/Q sky130_fd_sc_hd__dfxtp_4
X_22143_ _21564_/A _22139_/X _22314_/B _22142_/X VGND VGND VPWR VPWR _22144_/A sky130_fd_sc_hd__o22a_4
XFILLER_69_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24586__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22074_ _14487_/X _22074_/B _22073_/X VGND VGND VPWR VPWR _22074_/X sky130_fd_sc_hd__or3_4
XFILLER_114_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24515__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21025_ _20940_/X _20988_/X _21024_/Y VGND VGND VPWR VPWR _21025_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15583__A _11986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16274__B1 _22399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_HCLK_A clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15616__A3 _15501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14199__A _13934_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14824__B2 _24126_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11616__A _13665_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22976_ _16621_/A _22975_/X _22839_/X _24575_/Q _21694_/X VGND VGND VPWR VPWR _22976_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_28_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22362__A3 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24715_ _23664_/CLK _24715_/D HRESETn VGND VGND VPWR VPWR _14681_/A sky130_fd_sc_hd__dfrtp_4
X_21927_ _21158_/A _21927_/B VGND VGND VPWR VPWR _21927_/X sky130_fd_sc_hd__or2_4
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12660_ _12544_/Y _12657_/X VGND VGND VPWR VPWR _12660_/X sky130_fd_sc_hd__or2_4
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24646_ _24644_/CLK _15252_/X HRESETn VGND VGND VPWR VPWR _13753_/C sky130_fd_sc_hd__dfrtp_4
X_21858_ _21858_/A _21720_/B VGND VGND VPWR VPWR _21858_/X sky130_fd_sc_hd__and2_4
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ HWDATA[7] VGND VGND VPWR VPWR _13663_/A sky130_fd_sc_hd__buf_2
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ _20757_/X _20805_/X _20807_/X _20808_/Y VGND VGND VPWR VPWR _20809_/X sky130_fd_sc_hd__a211o_4
XFILLER_70_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17022__B _17022_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12552_/X _12591_/B _12591_/C _12590_/X VGND VGND VPWR VPWR _12591_/X sky130_fd_sc_hd__or4_4
XANTENNA__14772__A1_N _15045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24577_ _23353_/CLK _15454_/X HRESETn VGND VGND VPWR VPWR _15449_/A sky130_fd_sc_hd__dfrtp_4
X_21789_ _21764_/A _21784_/X _21786_/X _21787_/X _21788_/X VGND VGND VPWR VPWR _21789_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12447__A _12415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22863__B _23020_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ _20331_/A _14325_/X _24778_/Q _14327_/X VGND VGND VPWR VPWR _14330_/X sky130_fd_sc_hd__o22a_4
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ _11541_/X VGND VGND VPWR VPWR _11542_/X sky130_fd_sc_hd__buf_2
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23528_ _23537_/CLK _18894_/X VGND VGND VPWR VPWR _18893_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__21873__A2 _21082_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261_ _14259_/Y _14260_/X _14213_/X _14260_/X VGND VGND VPWR VPWR _24802_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23459_ _23457_/CLK _23459_/D VGND VGND VPWR VPWR _17828_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_137_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16000_ _15999_/Y _15922_/X _15709_/X _15922_/X VGND VGND VPWR VPWR _24361_/D sky130_fd_sc_hd__a2bb2o_4
X_13212_ _13244_/A _13212_/B VGND VGND VPWR VPWR _13212_/X sky130_fd_sc_hd__or2_4
X_14192_ _24824_/Q _14150_/X _14176_/X _11983_/A _14174_/Y VGND VGND VPWR VPWR _14192_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_87_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11574__B1 _11573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13143_ _13247_/A _13138_/X _13142_/X VGND VGND VPWR VPWR _13143_/X sky130_fd_sc_hd__or3_4
XANTENNA__17973__A _16231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25129_ _25130_/CLK _12212_/X HRESETn VGND VGND VPWR VPWR _25129_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_83_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12118__A2 _12117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21495__A _22148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13074_ _13271_/A VGND VGND VPWR VPWR _13207_/A sky130_fd_sc_hd__buf_2
X_17951_ _17887_/A _23415_/Q VGND VGND VPWR VPWR _17951_/X sky130_fd_sc_hd__or2_4
XFILLER_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24256__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12025_ _12015_/B VGND VGND VPWR VPWR _12025_/Y sky130_fd_sc_hd__inv_2
X_16902_ _16784_/Y _16902_/B VGND VGND VPWR VPWR _16903_/C sky130_fd_sc_hd__nand2_4
XFILLER_26_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17882_ _17914_/A _17880_/X _17882_/C VGND VGND VPWR VPWR _17883_/C sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_5_30_0_HCLK_A clkbuf_5_30_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12910__A _12921_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16265__B1 _16264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19621_ _23270_/Q VGND VGND VPWR VPWR _22087_/B sky130_fd_sc_hd__inv_2
X_16833_ _16833_/A VGND VGND VPWR VPWR _16834_/C sky130_fd_sc_hd__inv_2
XFILLER_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14815__A1 _24711_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16764_ _16757_/X _16759_/X _16762_/X _16764_/D VGND VGND VPWR VPWR _16764_/X sky130_fd_sc_hd__or4_4
X_19552_ _23294_/Q VGND VGND VPWR VPWR _22109_/B sky130_fd_sc_hd__inv_2
XANTENNA__22889__A1 _22195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13976_ _13973_/X _13975_/Y _24801_/Q _13973_/X VGND VGND VPWR VPWR _13976_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22889__B2 _22198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15715_ _24465_/Q VGND VGND VPWR VPWR _15717_/A sky130_fd_sc_hd__inv_2
X_18503_ _18503_/A _18503_/B VGND VGND VPWR VPWR _18503_/X sky130_fd_sc_hd__or2_4
XFILLER_74_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12927_ _12916_/B VGND VGND VPWR VPWR _12931_/B sky130_fd_sc_hd__inv_2
X_16695_ _16001_/Y _20778_/A _16001_/Y _20778_/A VGND VGND VPWR VPWR _16696_/D sky130_fd_sc_hd__a2bb2o_4
X_19483_ _19482_/Y _19480_/X _19366_/X _19480_/X VGND VGND VPWR VPWR _23320_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16736__A2_N _22853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_159_0_HCLK clkbuf_7_79_0_HCLK/X VGND VGND VPWR VPWR _24432_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__20540__A1_N _20419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15646_ _15461_/X _15641_/X _15635_/X _20739_/B _15645_/X VGND VGND VPWR VPWR _15646_/X
+ sky130_fd_sc_hd__a32o_4
X_18434_ _18358_/Y _18495_/B _18434_/C _18434_/D VGND VGND VPWR VPWR _18434_/X sky130_fd_sc_hd__or4_4
XANTENNA__23891__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12858_ _12858_/A VGND VGND VPWR VPWR _12858_/X sky130_fd_sc_hd__buf_2
XFILLER_62_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11809_ _11809_/A _11809_/B VGND VGND VPWR VPWR _11809_/X sky130_fd_sc_hd__and2_4
X_18365_ _23820_/Q VGND VGND VPWR VPWR _18535_/A sky130_fd_sc_hd__inv_2
XANTENNA__23820__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15577_ _15576_/X VGND VGND VPWR VPWR _15578_/B sky130_fd_sc_hd__buf_2
XFILLER_15_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12789_ _22258_/A _12787_/Y _12788_/Y _24455_/Q VGND VGND VPWR VPWR _12789_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12357__A _24472_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25044__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _23990_/Q VGND VGND VPWR VPWR _17325_/B sky130_fd_sc_hd__inv_2
X_14528_ _14528_/A VGND VGND VPWR VPWR _21007_/A sky130_fd_sc_hd__inv_2
X_18296_ _18290_/X _18296_/B _18296_/C VGND VGND VPWR VPWR _18296_/X sky130_fd_sc_hd__and3_4
XANTENNA__20574__A _20552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17247_ _17352_/A VGND VGND VPWR VPWR _17353_/A sky130_fd_sc_hd__inv_2
X_14459_ _24739_/Q VGND VGND VPWR VPWR _14542_/A sky130_fd_sc_hd__inv_2
XFILLER_70_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16293__A1_N _14936_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14572__A _14571_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16740__B2 _17614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17178_ _23674_/Q _20374_/A VGND VGND VPWR VPWR _17179_/B sky130_fd_sc_hd__or2_4
XFILLER_116_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22813__A1 _22931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16129_ _14197_/A _15822_/X VGND VGND VPWR VPWR _16129_/X sky130_fd_sc_hd__or2_4
XANTENNA__12109__A2 _24574_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16499__A _16499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13916__A _13908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19819_ _21957_/B _19814_/X _19818_/X _19814_/X VGND VGND VPWR VPWR _19819_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22592__A3 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23979__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22830_ _22826_/X _22830_/B _22830_/C _22829_/X VGND VGND VPWR VPWR _22830_/X sky130_fd_sc_hd__or4_4
XANTENNA__16271__A3 _15494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_55_0_HCLK clkbuf_7_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_55_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__20749__A _20818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23908__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22761_ _21972_/X _22760_/X _22634_/X _24525_/Q _21187_/X VGND VGND VPWR VPWR _22761_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_77_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14747__A _14747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24500_ _23949_/CLK _24500_/D HRESETn VGND VGND VPWR VPWR _24500_/Q sky130_fd_sc_hd__dfrtp_4
X_21712_ _22968_/A _21712_/B VGND VGND VPWR VPWR _21712_/Y sky130_fd_sc_hd__nand2_4
XFILLER_77_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11659__A2_N _21871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22692_ _24211_/Q _22580_/B VGND VGND VPWR VPWR _22692_/X sky130_fd_sc_hd__or2_4
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24431_ _24372_/CLK _15802_/X HRESETn VGND VGND VPWR VPWR _21269_/A sky130_fd_sc_hd__dfrtp_4
X_21643_ _18093_/A _20072_/Y _21644_/A _21181_/A VGND VGND VPWR VPWR _21643_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21304__B2 _21083_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24362_ _24412_/CLK _24362_/D HRESETn VGND VGND VPWR VPWR _24362_/Q sky130_fd_sc_hd__dfrtp_4
X_21574_ _24129_/Q _21553_/A _21292_/X _21573_/X VGND VGND VPWR VPWR _21574_/X sky130_fd_sc_hd__a211o_4
XANTENNA__20484__A _20511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23313_ _23313_/CLK _19502_/X VGND VGND VPWR VPWR _23313_/Q sky130_fd_sc_hd__dfxtp_4
X_20525_ _20524_/A _20524_/B _20524_/Y VGND VGND VPWR VPWR _20525_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_138_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15578__A _15414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24293_ _24590_/CLK _16209_/X HRESETn VGND VGND VPWR VPWR _24293_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24767__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20456_ _20456_/A VGND VGND VPWR VPWR _20456_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23244_ _23242_/CLK _19695_/X VGND VGND VPWR VPWR _19693_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__11556__B1 _11555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13098__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20387_ _15281_/Y _20367_/X _20357_/X _20386_/X VGND VGND VPWR VPWR _20388_/A sky130_fd_sc_hd__a211o_4
XFILLER_84_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23175_ _25106_/CLK _19881_/X VGND VGND VPWR VPWR _19880_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_49_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22126_ _22126_/A _21984_/X VGND VGND VPWR VPWR _22126_/X sky130_fd_sc_hd__or2_4
XFILLER_106_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22057_ _22064_/A _22057_/B VGND VGND VPWR VPWR _22057_/X sky130_fd_sc_hd__or2_4
XFILLER_88_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19433__B1 _19387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16202__A _16202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21008_ _21008_/A _21008_/B VGND VGND VPWR VPWR _21010_/B sky130_fd_sc_hd__or2_4
XANTENNA__13545__B _20554_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13830_ _13815_/A _13812_/X _13830_/C _13829_/X VGND VGND VPWR VPWR _13830_/X sky130_fd_sc_hd__or4_4
XFILLER_60_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23649__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13761_ _13761_/A _13761_/B _13716_/X _13782_/B VGND VGND VPWR VPWR _13762_/D sky130_fd_sc_hd__or4_4
XFILLER_55_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22959_ _21569_/A _22956_/X _22958_/X VGND VGND VPWR VPWR _22959_/X sky130_fd_sc_hd__and3_4
X_15500_ _15482_/X _15483_/X _15499_/X _24559_/Q _15495_/X VGND VGND VPWR VPWR _15500_/X
+ sky130_fd_sc_hd__a32o_4
X_12712_ _12565_/Y _12716_/B _12711_/Y VGND VGND VPWR VPWR _25056_/D sky130_fd_sc_hd__o21a_4
X_16480_ _16530_/A VGND VGND VPWR VPWR _16493_/A sky130_fd_sc_hd__buf_2
XFILLER_43_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13692_ _20402_/A _13687_/X _24920_/Q _13689_/X VGND VGND VPWR VPWR _13692_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22874__A _22997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15431_ HWDATA[0] VGND VGND VPWR VPWR _15431_/X sky130_fd_sc_hd__buf_2
X_12643_ _25058_/Q VGND VGND VPWR VPWR _12704_/A sky130_fd_sc_hd__inv_2
XFILLER_54_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24629_ _23676_/CLK _15280_/X HRESETn VGND VGND VPWR VPWR _24629_/Q sky130_fd_sc_hd__dfstp_4
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18150_ _23869_/Q VGND VGND VPWR VPWR _18242_/B sky130_fd_sc_hd__inv_2
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15362_ _15361_/Y _15359_/X _11573_/X _15359_/X VGND VGND VPWR VPWR _15362_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ _25044_/Q VGND VGND VPWR VPWR _12647_/C sky130_fd_sc_hd__inv_2
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17101_ _17101_/A _17101_/B _17100_/X VGND VGND VPWR VPWR _24048_/D sky130_fd_sc_hd__and3_4
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14313_ _23077_/Q _20179_/C _14311_/X _23617_/D _14312_/Y VGND VGND VPWR VPWR _24783_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11525_ HWDATA[29] VGND VGND VPWR VPWR _11525_/X sky130_fd_sc_hd__buf_2
X_18081_ _11737_/Y _18080_/Y VGND VGND VPWR VPWR _18081_/X sky130_fd_sc_hd__or2_4
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15293_ _24624_/Q _15245_/X _15243_/X VGND VGND VPWR VPWR _15293_/X sky130_fd_sc_hd__a21bo_4
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17032_ _17030_/Y _17161_/A _17160_/A _17032_/D VGND VGND VPWR VPWR _17035_/C sky130_fd_sc_hd__or4_4
XFILLER_32_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14244_ _13996_/Y _14243_/X _14213_/X _14243_/X VGND VGND VPWR VPWR _24810_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24437__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14175_ _14174_/Y VGND VGND VPWR VPWR _14175_/X sky130_fd_sc_hd__buf_2
X_13126_ _13073_/A _13122_/X _13125_/X VGND VGND VPWR VPWR _13126_/X sky130_fd_sc_hd__or3_4
X_18983_ _18981_/Y _18982_/X _18959_/X _18982_/X VGND VGND VPWR VPWR _18983_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22114__A _11532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24090__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13057_ _13057_/A VGND VGND VPWR VPWR _13057_/X sky130_fd_sc_hd__buf_2
X_17934_ _17934_/A _23512_/Q VGND VGND VPWR VPWR _17936_/B sky130_fd_sc_hd__or2_4
XFILLER_117_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22023__A2 _22007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16238__B1 _24286_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12008_ _12006_/Y _12002_/X _11636_/X _12007_/X VGND VGND VPWR VPWR _25140_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21953__A _21214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17865_ _17929_/A _17865_/B _17864_/X VGND VGND VPWR VPWR _17865_/X sky130_fd_sc_hd__and3_4
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17986__B1 _23922_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19604_ _19613_/A VGND VGND VPWR VPWR _19604_/X sky130_fd_sc_hd__buf_2
X_16816_ _24089_/Q VGND VGND VPWR VPWR _16816_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16253__A3 _15600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17796_ _17721_/A VGND VGND VPWR VPWR _17796_/X sky130_fd_sc_hd__buf_2
X_19535_ _22094_/B _19534_/X _11835_/X _19534_/X VGND VGND VPWR VPWR _19535_/X sky130_fd_sc_hd__a2bb2o_4
X_13959_ _13959_/A VGND VGND VPWR VPWR _23647_/D sky130_fd_sc_hd__buf_2
X_16747_ _16746_/X VGND VGND VPWR VPWR _16747_/Y sky130_fd_sc_hd__inv_2
X_16678_ _17725_/A VGND VGND VPWR VPWR _16678_/X sky130_fd_sc_hd__buf_2
X_19466_ _23326_/Q VGND VGND VPWR VPWR _19466_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16410__B1 _16153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18417_ _18363_/Y VGND VGND VPWR VPWR _18470_/A sky130_fd_sc_hd__buf_2
X_15629_ _12596_/Y _15628_/X _15393_/X _15628_/X VGND VGND VPWR VPWR _24507_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19397_ _19396_/Y VGND VGND VPWR VPWR _19397_/X sky130_fd_sc_hd__buf_2
XFILLER_37_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18348_ _16432_/Y _23829_/Q _16432_/Y _23829_/Q VGND VGND VPWR VPWR _18357_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18279_ _18279_/A _18282_/B VGND VGND VPWR VPWR _18279_/Y sky130_fd_sc_hd__nand2_4
X_20310_ _18615_/A _18614_/X VGND VGND VPWR VPWR _20310_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22008__B _21868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24860__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21290_ _21066_/B VGND VGND VPWR VPWR _22167_/A sky130_fd_sc_hd__buf_2
XANTENNA__11538__B1 _25218_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22798__B1 _20745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24178__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20241_ _20241_/A VGND VGND VPWR VPWR _20241_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19540__A2_N _19534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24107__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20172_ _20164_/B _20163_/C _20171_/B VGND VGND VPWR VPWR _20172_/X sky130_fd_sc_hd__o21a_4
XFILLER_103_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22024__A _20195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17118__A _24042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24980_ _24980_/CLK _24980_/D HRESETn VGND VGND VPWR VPWR _24980_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22959__A _21569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23931_ _24735_/CLK _23931_/D HRESETn VGND VGND VPWR VPWR _23931_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22970__B1 _11496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23862_ _23859_/CLK _23862_/D HRESETn VGND VGND VPWR VPWR _23862_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23742__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22813_ _22931_/A _22806_/X _22808_/X _22585_/X _22812_/Y VGND VGND VPWR VPWR _22813_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23793_ _23796_/CLK _20693_/Y HRESETn VGND VGND VPWR VPWR _12013_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_65_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22744_ _22722_/Y _22744_/B _22744_/C _22743_/X VGND VGND VPWR VPWR HRDATA[22] sky130_fd_sc_hd__or4_4
XFILLER_13_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14196__B _21072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_142_0_HCLK clkbuf_7_71_0_HCLK/X VGND VGND VPWR VPWR _23479_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22675_ _24309_/Q _22957_/B VGND VGND VPWR VPWR _22675_/X sky130_fd_sc_hd__and2_4
XANTENNA__16692__A _16692_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24948__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24414_ _24425_/CLK _15861_/X HRESETn VGND VGND VPWR VPWR _24414_/Q sky130_fd_sc_hd__dfrtp_4
X_21626_ _21626_/A _21624_/X _21625_/X VGND VGND VPWR VPWR _21626_/X sky130_fd_sc_hd__and3_4
XFILLER_16_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24345_ _24222_/CLK _16072_/X HRESETn VGND VGND VPWR VPWR _24345_/Q sky130_fd_sc_hd__dfrtp_4
X_21557_ _15278_/Y _21178_/A _24859_/Q _21400_/X VGND VGND VPWR VPWR _21557_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20508_ _20508_/A _20503_/Y VGND VGND VPWR VPWR _20508_/X sky130_fd_sc_hd__and2_4
XANTENNA__14715__B1 _14997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12290_ _12290_/A VGND VGND VPWR VPWR _25106_/D sky130_fd_sc_hd__inv_2
X_24276_ _24712_/CLK _24276_/D HRESETn VGND VGND VPWR VPWR _14900_/A sky130_fd_sc_hd__dfrtp_4
X_21488_ _17636_/X _21480_/X _21487_/X VGND VGND VPWR VPWR _21488_/X sky130_fd_sc_hd__or3_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24530__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23227_ _23246_/CLK _23227_/D VGND VGND VPWR VPWR _23227_/Q sky130_fd_sc_hd__dfxtp_4
X_20439_ _20438_/Y _20433_/Y _13505_/B VGND VGND VPWR VPWR _20439_/X sky130_fd_sc_hd__o21a_4
XFILLER_106_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16468__B1 _16211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23158_ _23179_/CLK _23158_/D VGND VGND VPWR VPWR _23158_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_121_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22109_ _20972_/A _22109_/B VGND VGND VPWR VPWR _22109_/X sky130_fd_sc_hd__or2_4
XFILLER_110_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15980_ _15977_/Y _15973_/X _15978_/X _15979_/X VGND VGND VPWR VPWR _15980_/X sky130_fd_sc_hd__a2bb2o_4
X_23089_ _23293_/CLK _23089_/D VGND VGND VPWR VPWR _23089_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20016__B2 _20015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14931_ _14931_/A _14924_/X _14927_/X _14931_/D VGND VGND VPWR VPWR _14931_/X sky130_fd_sc_hd__or4_4
XFILLER_103_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14862_ _14856_/X _14857_/X _14858_/X _14862_/D VGND VGND VPWR VPWR _14862_/X sky130_fd_sc_hd__or4_4
X_17650_ _23938_/Q VGND VGND VPWR VPWR _17651_/A sky130_fd_sc_hd__buf_2
XFILLER_90_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13813_ _13812_/X VGND VGND VPWR VPWR _13813_/Y sky130_fd_sc_hd__inv_2
X_16601_ _16601_/A VGND VGND VPWR VPWR _16601_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16640__B1 _16334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17581_ _17581_/A _17578_/X VGND VGND VPWR VPWR _17581_/X sky130_fd_sc_hd__or2_4
XFILLER_1_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14793_ _14786_/X _14788_/X _14789_/X _14792_/X VGND VGND VPWR VPWR _14794_/D sky130_fd_sc_hd__or4_4
XFILLER_75_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16532_ _16532_/A VGND VGND VPWR VPWR _16532_/Y sky130_fd_sc_hd__inv_2
X_19320_ _19318_/Y _19319_/X _19227_/X _19319_/X VGND VGND VPWR VPWR _23377_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13291__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13744_ _13745_/D _13739_/X _14074_/A VGND VGND VPWR VPWR _13744_/X sky130_fd_sc_hd__a21o_4
X_16463_ _16462_/Y _16460_/X _16376_/X _16460_/X VGND VGND VPWR VPWR _24195_/D sky130_fd_sc_hd__a2bb2o_4
X_19251_ _19238_/Y VGND VGND VPWR VPWR _19251_/X sky130_fd_sc_hd__buf_2
X_13675_ _13441_/Y _13649_/A _13645_/X _13649_/A VGND VGND VPWR VPWR _24925_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15414_ _15414_/A _21280_/A VGND VGND VPWR VPWR _16475_/B sky130_fd_sc_hd__or2_4
X_18202_ _23861_/Q VGND VGND VPWR VPWR _18202_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24689__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12626_ _12657_/A _24532_/Q _12657_/A _24532_/Q VGND VGND VPWR VPWR _12626_/X sky130_fd_sc_hd__a2bb2o_4
X_19182_ _19175_/A VGND VGND VPWR VPWR _19182_/X sky130_fd_sc_hd__buf_2
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16394_ _16393_/X VGND VGND VPWR VPWR _16401_/A sky130_fd_sc_hd__buf_2
XFILLER_31_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22109__A _20972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18133_ _16037_/Y _23876_/Q _16037_/Y _23876_/Q VGND VGND VPWR VPWR _18137_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24618__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15345_ _15353_/A VGND VGND VPWR VPWR _15345_/X sky130_fd_sc_hd__buf_2
X_12557_ _25063_/Q VGND VGND VPWR VPWR _12679_/C sky130_fd_sc_hd__inv_2
XANTENNA__22492__A2 _21882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19893__B1 _19825_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11508_ _11507_/X VGND VGND VPWR VPWR _16231_/A sky130_fd_sc_hd__buf_2
X_18064_ _23896_/Q VGND VGND VPWR VPWR _18064_/X sky130_fd_sc_hd__buf_2
XFILLER_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_4_0_HCLK_A clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15276_ _15285_/A VGND VGND VPWR VPWR _15276_/X sky130_fd_sc_hd__buf_2
X_12488_ _12373_/A _12487_/Y VGND VGND VPWR VPWR _12488_/X sky130_fd_sc_hd__or2_4
XFILLER_8_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20852__A _20852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17015_ _24317_/Q _17022_/B _16207_/Y _17027_/A VGND VGND VPWR VPWR _17017_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24271__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14227_ HWDATA[7] VGND VGND VPWR VPWR _16369_/A sky130_fd_sc_hd__buf_2
XANTENNA__19418__A _19417_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24200__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14158_ _12048_/B VGND VGND VPWR VPWR _14160_/B sky130_fd_sc_hd__inv_2
XFILLER_4_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13109_ _13016_/A VGND VGND VPWR VPWR _13110_/A sky130_fd_sc_hd__buf_2
XFILLER_113_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14089_ _14088_/Y _14084_/X _13635_/X _14084_/X VGND VGND VPWR VPWR _24858_/D sky130_fd_sc_hd__a2bb2o_4
X_18966_ _13041_/B VGND VGND VPWR VPWR _18966_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17917_ _17853_/A _23424_/Q VGND VGND VPWR VPWR _17918_/C sky130_fd_sc_hd__or2_4
X_18897_ _17682_/B VGND VGND VPWR VPWR _18897_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22498__B _22497_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17848_ _17944_/A _17848_/B VGND VGND VPWR VPWR _17848_/X sky130_fd_sc_hd__or2_4
XFILLER_39_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15434__A1 _15430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16631__B1 _11536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17779_ _17817_/A _19174_/A VGND VGND VPWR VPWR _17780_/C sky130_fd_sc_hd__or2_4
XANTENNA__13445__B1 _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19518_ _19518_/A VGND VGND VPWR VPWR _21676_/B sky130_fd_sc_hd__inv_2
X_20790_ _24393_/Q _20826_/A _20737_/A _15637_/X VGND VGND VPWR VPWR _20790_/X sky130_fd_sc_hd__o22a_4
X_19449_ _19440_/Y VGND VGND VPWR VPWR _19449_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_215_0_HCLK clkbuf_8_215_0_HCLK/A VGND VGND VPWR VPWR _23826_/CLK sky130_fd_sc_hd__clkbuf_1
X_22460_ _21047_/A VGND VGND VPWR VPWR _22460_/X sky130_fd_sc_hd__buf_2
XANTENNA__24359__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21411_ _24363_/Q _21043_/X VGND VGND VPWR VPWR _21411_/X sky130_fd_sc_hd__or2_4
X_22391_ _24480_/Q _22999_/B VGND VGND VPWR VPWR _22391_/X sky130_fd_sc_hd__or2_4
XFILLER_124_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24130_ _24101_/CLK _16612_/X HRESETn VGND VGND VPWR VPWR _24130_/Q sky130_fd_sc_hd__dfrtp_4
X_21342_ _21342_/A _21342_/B VGND VGND VPWR VPWR _21342_/X sky130_fd_sc_hd__or2_4
XFILLER_15_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24061_ _24618_/CLK _16953_/X HRESETn VGND VGND VPWR VPWR _24061_/Q sky130_fd_sc_hd__dfrtp_4
X_21273_ _21273_/A VGND VGND VPWR VPWR _23023_/A sky130_fd_sc_hd__buf_2
X_23012_ _23012_/A _23004_/A VGND VGND VPWR VPWR _23012_/X sky130_fd_sc_hd__and2_4
X_20224_ _20266_/A _20224_/B _20266_/C VGND VGND VPWR VPWR _20224_/X sky130_fd_sc_hd__or3_4
XFILLER_131_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20155_ _23761_/D _20155_/B VGND VGND VPWR VPWR _20155_/X sky130_fd_sc_hd__or2_4
XFILLER_89_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23994__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23923__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20086_ _23097_/Q VGND VGND VPWR VPWR _20086_/Y sky130_fd_sc_hd__inv_2
X_24963_ _24980_/CLK _24963_/D HRESETn VGND VGND VPWR VPWR _20881_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25147__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12430__D _12417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23914_ _23908_/CLK _23914_/D HRESETn VGND VGND VPWR VPWR _23914_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24894_ _23624_/CLK _24894_/D HRESETn VGND VGND VPWR VPWR _13924_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_79_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23845_ _23845_/CLK _23845_/D HRESETn VGND VGND VPWR VPWR _23845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_25_0_HCLK clkbuf_6_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11624__A HWDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11790_ _11809_/A VGND VGND VPWR VPWR _11815_/C sky130_fd_sc_hd__buf_2
XFILLER_60_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23776_ _23668_/CLK _23776_/D HRESETn VGND VGND VPWR VPWR _20164_/B sky130_fd_sc_hd__dfrtp_4
X_20988_ _17631_/Y _20955_/X _20969_/X _20981_/X _20987_/X VGND VGND VPWR VPWR _20988_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__11998__B1 _11616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22727_ _16583_/Y _21544_/X _14960_/Y _22312_/B VGND VGND VPWR VPWR _22727_/X sky130_fd_sc_hd__o22a_4
XFILLER_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24782__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13460_ _24620_/Q _24619_/Q _22510_/B VGND VGND VPWR VPWR _13460_/X sky130_fd_sc_hd__or3_4
XFILLER_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22658_ _22656_/Y _22610_/X _23746_/Q _22657_/X VGND VGND VPWR VPWR _22658_/X sky130_fd_sc_hd__a2bb2o_4
X_12411_ _12411_/A _12411_/B _12410_/Y _12385_/Y VGND VGND VPWR VPWR _12411_/X sky130_fd_sc_hd__or4_4
XANTENNA__24711__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21609_ _21625_/A _21609_/B VGND VGND VPWR VPWR _21609_/X sky130_fd_sc_hd__or2_4
XFILLER_107_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13391_ _13391_/A _13391_/B VGND VGND VPWR VPWR _13391_/X sky130_fd_sc_hd__and2_4
XFILLER_16_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22589_ _22588_/X VGND VGND VPWR VPWR _22589_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24029__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15130_ _15130_/A VGND VGND VPWR VPWR _15130_/Y sky130_fd_sc_hd__inv_2
X_12342_ _24496_/Q VGND VGND VPWR VPWR _12342_/Y sky130_fd_sc_hd__inv_2
X_24328_ _23852_/CLK _24328_/D HRESETn VGND VGND VPWR VPWR _24328_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_103_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15061_ _14873_/D _15061_/B VGND VGND VPWR VPWR _15064_/B sky130_fd_sc_hd__or2_4
X_12273_ _12178_/C _12276_/B _12195_/X VGND VGND VPWR VPWR _12273_/Y sky130_fd_sc_hd__a21oi_4
X_24259_ _24259_/CLK _24259_/D HRESETn VGND VGND VPWR VPWR _24259_/Q sky130_fd_sc_hd__dfrtp_4
X_14012_ _20232_/A VGND VGND VPWR VPWR _14012_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18820_ _18819_/Y _18814_/X _18795_/X _18814_/X VGND VGND VPWR VPWR _18820_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18751_ _23577_/Q VGND VGND VPWR VPWR _18751_/Y sky130_fd_sc_hd__inv_2
X_15963_ _22458_/A VGND VGND VPWR VPWR _15963_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_107_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_215_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13675__B1 _13645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17702_ _17702_/A _17702_/B _17701_/X VGND VGND VPWR VPWR _17702_/X sky130_fd_sc_hd__and3_4
X_14914_ _24674_/Q _24279_/Q _15138_/B _14913_/Y VGND VGND VPWR VPWR _14918_/C sky130_fd_sc_hd__o22a_4
X_15894_ _16373_/A VGND VGND VPWR VPWR _15894_/X sky130_fd_sc_hd__buf_2
X_18682_ _18682_/A VGND VGND VPWR VPWR _18682_/X sky130_fd_sc_hd__buf_2
XANTENNA__16630__A1_N _14740_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16613__B1 _16546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17633_ _23941_/Q _17632_/A _17631_/Y _17632_/Y VGND VGND VPWR VPWR _17634_/A sky130_fd_sc_hd__o22a_4
XANTENNA__22903__A2_N _20926_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14845_ _15067_/C _16608_/A _15067_/C _16608_/A VGND VGND VPWR VPWR _14845_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11534__A _15916_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19701__A _19688_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14776_ _24686_/Q VGND VGND VPWR VPWR _15059_/A sky130_fd_sc_hd__inv_2
X_17564_ _17547_/X _17564_/B _17563_/Y VGND VGND VPWR VPWR _23960_/D sky130_fd_sc_hd__and3_4
X_11988_ _21564_/A VGND VGND VPWR VPWR _15271_/A sky130_fd_sc_hd__buf_2
XANTENNA__22162__A1 _24510_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19303_ _19303_/A _18075_/X _18068_/X _18064_/X VGND VGND VPWR VPWR _19304_/A sky130_fd_sc_hd__or4_4
X_13727_ _13726_/X VGND VGND VPWR VPWR _13732_/A sky130_fd_sc_hd__inv_2
X_16515_ _24174_/Q VGND VGND VPWR VPWR _16515_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17495_ _22473_/A VGND VGND VPWR VPWR _17497_/A sky130_fd_sc_hd__inv_2
XFILLER_17_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19234_ _23406_/Q VGND VGND VPWR VPWR _19234_/Y sky130_fd_sc_hd__inv_2
X_13658_ _15788_/A VGND VGND VPWR VPWR _13658_/X sky130_fd_sc_hd__buf_2
X_16446_ _16452_/A VGND VGND VPWR VPWR _16446_/X sky130_fd_sc_hd__buf_2
XANTENNA__24452__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12609_ _12609_/A VGND VGND VPWR VPWR _12609_/Y sky130_fd_sc_hd__inv_2
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16377_ _16375_/Y _16372_/X _16376_/X _16372_/X VGND VGND VPWR VPWR _16377_/X sky130_fd_sc_hd__a2bb2o_4
X_19165_ _19164_/Y _19160_/X _19120_/X _19153_/A VGND VGND VPWR VPWR _19165_/X sky130_fd_sc_hd__a2bb2o_4
X_13589_ _11679_/Y _13561_/B VGND VGND VPWR VPWR _13589_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_45_0_HCLK clkbuf_8_45_0_HCLK/A VGND VGND VPWR VPWR _24998_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15328_ _15324_/Y _15327_/X _11522_/X _15327_/X VGND VGND VPWR VPWR _24614_/D sky130_fd_sc_hd__a2bb2o_4
X_18116_ _21898_/A _18113_/X _23883_/Q _18113_/X VGND VGND VPWR VPWR _18116_/X sky130_fd_sc_hd__a2bb2o_4
X_19096_ _19094_/Y _19092_/X _19095_/X _19092_/X VGND VGND VPWR VPWR _23456_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15259_ _13726_/X _15247_/X _15256_/X _13716_/D _15254_/X VGND VGND VPWR VPWR _15259_/X
+ sky130_fd_sc_hd__a32o_4
X_18047_ _23940_/Q VGND VGND VPWR VPWR _18047_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22475__A1_N _12489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19998_ _23131_/Q VGND VGND VPWR VPWR _19998_/Y sky130_fd_sc_hd__inv_2
X_18949_ _18949_/A VGND VGND VPWR VPWR _18949_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13666__B1 _13665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21960_ _21777_/A _21960_/B VGND VGND VPWR VPWR _21960_/X sky130_fd_sc_hd__or2_4
XANTENNA__22659__D _22658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16604__B1 _16279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20911_ _21357_/A VGND VGND VPWR VPWR _20911_/X sky130_fd_sc_hd__buf_2
XFILLER_66_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21891_ _24822_/Q _22024_/B VGND VGND VPWR VPWR _21891_/X sky130_fd_sc_hd__and2_4
XFILLER_54_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14938__A2_N _14936_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23630_ _23641_/CLK _23630_/D HRESETn VGND VGND VPWR VPWR _18608_/B sky130_fd_sc_hd__dfrtp_4
X_20842_ _16043_/A _20842_/B _20842_/C VGND VGND VPWR VPWR _21079_/B sky130_fd_sc_hd__or3_4
XANTENNA__21860__B _21860_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20757__A _20757_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23561_ _23586_/CLK _18799_/X VGND VGND VPWR VPWR _23561_/Q sky130_fd_sc_hd__dfxtp_4
X_20773_ _11514_/X VGND VGND VPWR VPWR _21990_/A sky130_fd_sc_hd__inv_2
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14755__A _24098_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22512_ _22512_/A _22997_/A VGND VGND VPWR VPWR _22832_/C sky130_fd_sc_hd__or2_4
XFILLER_52_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23492_ _23493_/CLK _18997_/X VGND VGND VPWR VPWR _23492_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22972__A _24459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24193__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22443_ _22443_/A VGND VGND VPWR VPWR _22456_/B sky130_fd_sc_hd__inv_2
XANTENNA__15591__B1 _11525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19857__B1 _19835_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24122__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21588__A _11952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25162_ _24623_/CLK _11925_/X HRESETn VGND VGND VPWR VPWR _11923_/A sky130_fd_sc_hd__dfrtp_4
X_22374_ _22129_/X _22373_/X _21994_/X _24557_/Q _21995_/X VGND VGND VPWR VPWR _22374_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_11_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24113_ _24113_/CLK _16641_/X HRESETn VGND VGND VPWR VPWR _24113_/Q sky130_fd_sc_hd__dfrtp_4
X_21325_ _21348_/A _21325_/B VGND VGND VPWR VPWR _21325_/X sky130_fd_sc_hd__or2_4
XANTENNA__15343__B1 _11552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25093_ _25097_/CLK _12460_/X HRESETn VGND VGND VPWR VPWR _25093_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24044_ _24308_/CLK _17113_/X HRESETn VGND VGND VPWR VPWR _16992_/A sky130_fd_sc_hd__dfrtp_4
X_21256_ _20782_/A VGND VGND VPWR VPWR _21256_/X sky130_fd_sc_hd__buf_2
X_20207_ _20200_/Y _14102_/X _20212_/D _20206_/X VGND VGND VPWR VPWR _20207_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11619__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21187_ _22198_/A VGND VGND VPWR VPWR _21187_/X sky130_fd_sc_hd__buf_2
XANTENNA__13537__C _13537_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15646__A1 _15461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20138_ _23075_/Q VGND VGND VPWR VPWR _20138_/Y sky130_fd_sc_hd__inv_2
X_12960_ _12833_/X _12955_/B _12922_/X _12957_/B VGND VGND VPWR VPWR _12961_/A sky130_fd_sc_hd__a211o_4
X_20069_ _20069_/A VGND VGND VPWR VPWR _20070_/A sky130_fd_sc_hd__inv_2
X_24946_ _24851_/CLK _13621_/X HRESETn VGND VGND VPWR VPWR _24946_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18596__B1 _24249_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11911_ _11909_/X VGND VGND VPWR VPWR _11911_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12891_ _12921_/A _12889_/X _12891_/C VGND VGND VPWR VPWR _25036_/D sky130_fd_sc_hd__and3_4
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24877_ _24879_/CLK _14033_/X HRESETn VGND VGND VPWR VPWR _20209_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14630_ _14630_/A _14630_/B _14608_/Y VGND VGND VPWR VPWR _14631_/B sky130_fd_sc_hd__and3_4
XANTENNA__24963__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11842_ _11842_/A VGND VGND VPWR VPWR _19607_/A sky130_fd_sc_hd__buf_2
XANTENNA__18119__A1_N _18117_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23828_ _23828_/CLK _23828_/D HRESETn VGND VGND VPWR VPWR _18430_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14082__B1 _13665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14561_ _14561_/A _14560_/Y VGND VGND VPWR VPWR _14561_/X sky130_fd_sc_hd__or2_4
X_11773_ _11809_/A _11771_/Y _11773_/C VGND VGND VPWR VPWR _11795_/B sky130_fd_sc_hd__or3_4
X_23759_ _24112_/CLK _23759_/D HRESETn VGND VGND VPWR VPWR _23759_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13512_ _23720_/Q _20524_/A _13512_/C _20524_/B VGND VGND VPWR VPWR _13512_/X sky130_fd_sc_hd__or4_4
X_16300_ _16300_/A VGND VGND VPWR VPWR _22230_/A sky130_fd_sc_hd__buf_2
XANTENNA__17041__A _17041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17280_ _11572_/Y _17270_/A _25211_/Q _17246_/Y VGND VGND VPWR VPWR _17280_/X sky130_fd_sc_hd__a2bb2o_4
X_14492_ _14488_/X _14491_/X _14488_/X _14491_/X VGND VGND VPWR VPWR _14497_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16231_ _16231_/A _22017_/A VGND VGND VPWR VPWR _16235_/B sky130_fd_sc_hd__or2_4
X_13443_ _13441_/Y _14424_/B _13441_/Y _14424_/B VGND VGND VPWR VPWR _13443_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11801__B RsRx_S1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_4_0_HCLK clkbuf_8_5_0_HCLK/A VGND VGND VPWR VPWR _23242_/CLK sky130_fd_sc_hd__clkbuf_1
X_16162_ _16162_/A VGND VGND VPWR VPWR _16162_/Y sky130_fd_sc_hd__inv_2
X_13374_ _24980_/Q VGND VGND VPWR VPWR _13374_/Y sky130_fd_sc_hd__inv_2
X_15113_ _15108_/X _15110_/X _15112_/X VGND VGND VPWR VPWR _15187_/B sky130_fd_sc_hd__or3_4
X_12325_ _25088_/Q VGND VGND VPWR VPWR _12412_/A sky130_fd_sc_hd__inv_2
X_16093_ _16093_/A VGND VGND VPWR VPWR _16093_/X sky130_fd_sc_hd__buf_2
XFILLER_126_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15334__B1 _15332_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12913__A _12922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15044_ _15044_/A _15044_/B VGND VGND VPWR VPWR _15046_/B sky130_fd_sc_hd__or2_4
X_19921_ _21229_/B _19918_/X _19835_/X _19918_/X VGND VGND VPWR VPWR _23160_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12256_ _12186_/B _12256_/B VGND VGND VPWR VPWR _12257_/B sky130_fd_sc_hd__or2_4
XANTENNA__23845__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25069__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11529__A _11529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19852_ _21509_/B _19847_/X _19828_/X _19847_/X VGND VGND VPWR VPWR _23186_/D sky130_fd_sc_hd__a2bb2o_4
X_12187_ _12189_/B VGND VGND VPWR VPWR _12188_/B sky130_fd_sc_hd__inv_2
XFILLER_29_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18803_ _18800_/Y _18798_/X _18802_/X _18798_/X VGND VGND VPWR VPWR _23560_/D sky130_fd_sc_hd__a2bb2o_4
X_19783_ _19783_/A VGND VGND VPWR VPWR _19783_/Y sky130_fd_sc_hd__inv_2
X_16995_ _24032_/Q VGND VGND VPWR VPWR _17134_/A sky130_fd_sc_hd__inv_2
XFILLER_84_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22122__A _22121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18734_ _19946_/A _19123_/D _19946_/C _18734_/D VGND VGND VPWR VPWR _18734_/X sky130_fd_sc_hd__or4_4
X_15946_ _15945_/Y _15941_/X _15765_/X _15941_/X VGND VGND VPWR VPWR _24382_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21961__A _21229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18665_ _11755_/Y _11729_/X _18065_/C VGND VGND VPWR VPWR _18666_/C sky130_fd_sc_hd__or3_4
XFILLER_48_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15877_ _24407_/Q VGND VGND VPWR VPWR _15877_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17616_ _17487_/Y _17615_/X _16748_/X VGND VGND VPWR VPWR _17616_/Y sky130_fd_sc_hd__a21oi_4
X_14828_ _24695_/Q _24138_/Q _15019_/A _14827_/Y VGND VGND VPWR VPWR _14828_/X sky130_fd_sc_hd__o22a_4
X_18596_ _24243_/Q _18491_/A _24249_/Q _18462_/A VGND VGND VPWR VPWR _18596_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18339__B1 _16445_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22135__B2 _22121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24633__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17547_ _17619_/A VGND VGND VPWR VPWR _17547_/X sky130_fd_sc_hd__buf_2
XANTENNA__20146__B1 _15522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14759_ _14759_/A VGND VGND VPWR VPWR _14759_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17478_ _22979_/A VGND VGND VPWR VPWR _17478_/Y sky130_fd_sc_hd__inv_2
X_19217_ _23412_/Q VGND VGND VPWR VPWR _21746_/A sky130_fd_sc_hd__inv_2
X_16429_ _16428_/Y _16426_/X _16264_/X _16426_/X VGND VGND VPWR VPWR _16429_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12095__A _24564_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19148_ _23437_/Q VGND VGND VPWR VPWR _19148_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14128__A1 MSO_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14128__B2 _14122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19079_ _19078_/Y VGND VGND VPWR VPWR _19079_/X sky130_fd_sc_hd__buf_2
XFILLER_121_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21110_ _21280_/A VGND VGND VPWR VPWR _22279_/A sky130_fd_sc_hd__buf_2
X_22090_ _18048_/X _22086_/X _22089_/X VGND VGND VPWR VPWR _22090_/X sky130_fd_sc_hd__or3_4
X_21041_ _20751_/X VGND VGND VPWR VPWR _21042_/A sky130_fd_sc_hd__buf_2
XFILLER_82_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24800_ _24811_/CLK _14265_/X HRESETn VGND VGND VPWR VPWR _24800_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_68_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22992_ _16477_/Y _22992_/B VGND VGND VPWR VPWR _22992_/X sky130_fd_sc_hd__and2_4
XANTENNA__12311__B1 _12451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21871__A _21871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24731_ _23586_/CLK _24731_/D HRESETn VGND VGND VPWR VPWR _18873_/B sky130_fd_sc_hd__dfrtp_4
X_21943_ _21371_/A _21943_/B VGND VGND VPWR VPWR _21943_/X sky130_fd_sc_hd__or2_4
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20924__A2 _20923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_7_0_HCLK_A clkbuf_5_6_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21590__B _21590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24662_ _24662_/CLK _24662_/D HRESETn VGND VGND VPWR VPWR _24662_/Q sky130_fd_sc_hd__dfrtp_4
X_21874_ _21192_/X _21871_/X _21873_/X VGND VGND VPWR VPWR _21874_/X sky130_fd_sc_hd__and3_4
XFILLER_43_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15800__A1 _15799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15800__B2 _15746_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24374__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ _23489_/CLK _18648_/X VGND VGND VPWR VPWR _23613_/Q sky130_fd_sc_hd__dfxtp_4
X_20825_ _21097_/B VGND VGND VPWR VPWR _21716_/B sky130_fd_sc_hd__buf_2
XANTENNA__20137__B1 _17993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24593_ _23734_/CLK _24593_/D HRESETn VGND VGND VPWR VPWR _24593_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17002__B1 _24310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24303__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21885__B1 _21883_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23544_ _23479_/CLK _23544_/D VGND VGND VPWR VPWR _23544_/Q sky130_fd_sc_hd__dfxtp_4
X_20756_ _22036_/A VGND VGND VPWR VPWR _20757_/A sky130_fd_sc_hd__buf_2
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18750__B1 _18679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17796__A _17721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23475_ _23471_/CLK _19045_/X VGND VGND VPWR VPWR _23475_/Q sky130_fd_sc_hd__dfxtp_4
X_20687_ _11891_/A _20688_/B VGND VGND VPWR VPWR _23784_/D sky130_fd_sc_hd__and2_4
XFILLER_126_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25214_ _25214_/CLK _11553_/X HRESETn VGND VGND VPWR VPWR _25214_/Q sky130_fd_sc_hd__dfrtp_4
X_22426_ _24559_/Q _20799_/X _20801_/X _22425_/X VGND VGND VPWR VPWR _22426_/X sky130_fd_sc_hd__a211o_4
XFILLER_104_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22207__A _16041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25145_ _24984_/CLK _11996_/X HRESETn VGND VGND VPWR VPWR _25145_/Q sky130_fd_sc_hd__dfrtp_4
X_22357_ _20917_/X _22355_/X _20902_/X _22356_/Y VGND VGND VPWR VPWR _22357_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_8_91_0_HCLK clkbuf_8_91_0_HCLK/A VGND VGND VPWR VPWR _24870_/CLK sky130_fd_sc_hd__clkbuf_1
X_12110_ _12110_/A VGND VGND VPWR VPWR _12176_/A sky130_fd_sc_hd__inv_2
X_21308_ _21447_/A VGND VGND VPWR VPWR _21308_/X sky130_fd_sc_hd__buf_2
X_13090_ _11751_/X VGND VGND VPWR VPWR _13090_/X sky130_fd_sc_hd__buf_2
X_25076_ _25090_/CLK _12523_/X HRESETn VGND VGND VPWR VPWR _25076_/Q sky130_fd_sc_hd__dfrtp_4
X_22288_ _22335_/A VGND VGND VPWR VPWR _22349_/B sky130_fd_sc_hd__buf_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25162__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12041_ _12041_/A VGND VGND VPWR VPWR _12041_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24027_ _24289_/CLK _24027_/D HRESETn VGND VGND VPWR VPWR _17031_/A sky130_fd_sc_hd__dfrtp_4
X_21239_ _21392_/A _19878_/Y VGND VGND VPWR VPWR _21241_/B sky130_fd_sc_hd__or2_4
XFILLER_46_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23683__D sda_i_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15800_ _15799_/X _15582_/A _15706_/X _24432_/Q _15746_/A VGND VGND VPWR VPWR _15800_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_63_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17036__A _24040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13992_ _13925_/A _13925_/B _13925_/C _13950_/A VGND VGND VPWR VPWR _13992_/X sky130_fd_sc_hd__or4_4
X_16780_ _16780_/A VGND VGND VPWR VPWR _16780_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21781__A _21383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12943_ _12796_/Y _12947_/A _12943_/C _12943_/D VGND VGND VPWR VPWR _12943_/X sky130_fd_sc_hd__or4_4
X_15731_ _15717_/A _15717_/B _15730_/X VGND VGND VPWR VPWR _15731_/X sky130_fd_sc_hd__o21a_4
XFILLER_111_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24929_ _24937_/CLK _24929_/D HRESETn VGND VGND VPWR VPWR _24929_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18450_ _18440_/A _18447_/X _18442_/B _18449_/X VGND VGND VPWR VPWR _18451_/A sky130_fd_sc_hd__a211o_4
X_12874_ _12858_/A _12818_/Y _12999_/A _12793_/Y VGND VGND VPWR VPWR _12878_/C sky130_fd_sc_hd__or4_4
X_15662_ _15658_/X _15647_/X _15320_/X _24498_/Q _15661_/X VGND VGND VPWR VPWR _24498_/D
+ sky130_fd_sc_hd__a32o_4
X_17401_ _17400_/X VGND VGND VPWR VPWR _17401_/Y sky130_fd_sc_hd__inv_2
X_11825_ _11776_/B _11823_/Y _11824_/Y VGND VGND VPWR VPWR _11825_/X sky130_fd_sc_hd__o21a_4
X_14613_ _24725_/Q _14612_/X _24726_/Q VGND VGND VPWR VPWR _14614_/B sky130_fd_sc_hd__or3_4
XFILLER_57_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15593_ _15593_/A VGND VGND VPWR VPWR _15593_/X sky130_fd_sc_hd__buf_2
X_18381_ _23814_/Q VGND VGND VPWR VPWR _18551_/A sky130_fd_sc_hd__inv_2
XFILLER_61_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20128__B1 _19963_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12908__A _22900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24044__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14544_/A _14543_/X _14493_/A _19779_/B VGND VGND VPWR VPWR _19813_/A sky130_fd_sc_hd__or4_4
X_17332_ _17237_/A _17331_/Y VGND VGND VPWR VPWR _17332_/X sky130_fd_sc_hd__or2_4
XPHY_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _23894_/Q VGND VGND VPWR VPWR _18075_/A sky130_fd_sc_hd__inv_2
XPHY_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18741__B1 _18740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14475_ _14429_/X _14437_/X _14466_/X _14474_/X VGND VGND VPWR VPWR _14475_/X sky130_fd_sc_hd__or4_4
X_17263_ _25199_/Q _23987_/Q _11603_/Y _17262_/Y VGND VGND VPWR VPWR _17263_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11687_ _11687_/A VGND VGND VPWR VPWR _11687_/Y sky130_fd_sc_hd__inv_2
XPHY_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19002_ _19002_/A VGND VGND VPWR VPWR _19002_/Y sky130_fd_sc_hd__inv_2
X_13426_ _22449_/A _24767_/Q _22449_/A _24767_/Q VGND VGND VPWR VPWR _13427_/D sky130_fd_sc_hd__a2bb2o_4
X_16214_ _16213_/Y _16208_/X _15801_/X _16208_/X VGND VGND VPWR VPWR _24291_/D sky130_fd_sc_hd__a2bb2o_4
X_17194_ _17170_/Y _17184_/Y _23682_/Q _20723_/B _17187_/X VGND VGND VPWR VPWR _24021_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_127_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19297__B2 _19296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22117__A _24367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16145_ _16165_/A VGND VGND VPWR VPWR _16145_/X sky130_fd_sc_hd__buf_2
X_13357_ _11503_/A VGND VGND VPWR VPWR _13357_/X sky130_fd_sc_hd__buf_2
XANTENNA__15307__B1 HADDR[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12308_ _25097_/Q VGND VGND VPWR VPWR _12417_/A sky130_fd_sc_hd__inv_2
XFILLER_115_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16076_ _16071_/A VGND VGND VPWR VPWR _16076_/X sky130_fd_sc_hd__buf_2
XFILLER_5_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_119_0_HCLK clkbuf_7_59_0_HCLK/X VGND VGND VPWR VPWR _24643_/CLK sky130_fd_sc_hd__clkbuf_1
X_13288_ _11710_/X _13272_/X _13287_/X _24998_/Q _11708_/X VGND VGND VPWR VPWR _13288_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_5_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15027_ _14984_/A VGND VGND VPWR VPWR _15027_/X sky130_fd_sc_hd__buf_2
X_19904_ _14548_/X _14543_/X _14493_/A _19904_/D VGND VGND VPWR VPWR _19904_/X sky130_fd_sc_hd__or4_4
X_12239_ _12174_/A _12174_/B _12083_/X _12252_/B VGND VGND VPWR VPWR _12245_/B sky130_fd_sc_hd__or4_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22151__A2_N _20940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19835_ _19835_/A VGND VGND VPWR VPWR _19835_/X sky130_fd_sc_hd__buf_2
XANTENNA__23627__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24885__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19766_ _21812_/B _19760_/X _19717_/X _19765_/X VGND VGND VPWR VPWR _19766_/X sky130_fd_sc_hd__a2bb2o_4
X_16978_ _24313_/Q _24051_/Q _16157_/Y _17026_/B VGND VGND VPWR VPWR _16978_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14294__B1 _14236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22787__A _20820_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18717_ _18716_/Y _14594_/X _17202_/X _14594_/X VGND VGND VPWR VPWR _18717_/X sky130_fd_sc_hd__a2bb2o_4
X_15929_ _15928_/X VGND VGND VPWR VPWR _15929_/X sky130_fd_sc_hd__buf_2
X_19697_ _19696_/Y _19694_/X _19607_/X _19694_/X VGND VGND VPWR VPWR _19697_/X sky130_fd_sc_hd__a2bb2o_4
X_18648_ _21949_/B _18645_/X _15545_/X _18645_/X VGND VGND VPWR VPWR _18648_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18980__B1 _18932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18579_ _16310_/A _23843_/Q _16310_/Y _18440_/A VGND VGND VPWR VPWR _18579_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15794__B1 _15390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20610_ _20606_/X VGND VGND VPWR VPWR _20610_/Y sky130_fd_sc_hd__inv_2
X_21590_ _16378_/Y _21590_/B VGND VGND VPWR VPWR _21592_/B sky130_fd_sc_hd__or2_4
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20541_ _20542_/A VGND VGND VPWR VPWR _20541_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12618__A2_N _24528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20754__B _23025_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23767__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23260_ _23258_/CLK _19653_/X VGND VGND VPWR VPWR _19651_/A sky130_fd_sc_hd__dfxtp_4
X_20472_ _13508_/D VGND VGND VPWR VPWR _20472_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22211_ _16532_/Y _15572_/A VGND VGND VPWR VPWR _22211_/X sky130_fd_sc_hd__and2_4
Xclkbuf_7_15_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_106_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23191_ _25106_/CLK _23191_/D VGND VGND VPWR VPWR _23191_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_78_0_HCLK clkbuf_7_78_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_78_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22142_ _21707_/B _22140_/X _11954_/X _22141_/X VGND VGND VPWR VPWR _22142_/X sky130_fd_sc_hd__o22a_4
XFILLER_134_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20770__A _20750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15864__A _24412_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22044__B1 _23917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22073_ _21764_/A _22071_/X _22073_/C VGND VGND VPWR VPWR _22073_/X sky130_fd_sc_hd__and3_4
XFILLER_0_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18240__A _18263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21398__A2 _14016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21024_ _21024_/A VGND VGND VPWR VPWR _21024_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15583__B _15741_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14285__B1 _14218_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14199__B _14199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24555__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18015__A2 _16228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22975_ _22975_/A _23008_/B VGND VGND VPWR VPWR _22975_/X sky130_fd_sc_hd__or2_4
XFILLER_56_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17223__B1 _16556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20929__B _22488_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21926_ _21346_/A _21924_/X _21925_/X VGND VGND VPWR VPWR _21926_/X sky130_fd_sc_hd__and3_4
XFILLER_76_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24714_ _24674_/CLK _14865_/Y HRESETn VGND VGND VPWR VPWR pwm_S6 sky130_fd_sc_hd__dfrtp_4
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18971__B1 _18901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24645_ _24643_/CLK _15253_/X HRESETn VGND VGND VPWR VPWR _13718_/B sky130_fd_sc_hd__dfrtp_4
X_21857_ _21857_/A _21745_/X _21857_/C _21856_/X VGND VGND VPWR VPWR HRDATA[5] sky130_fd_sc_hd__or4_4
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11599_/A VGND VGND VPWR VPWR _11610_/X sky130_fd_sc_hd__buf_2
XFILLER_58_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _20808_/A _13618_/A VGND VGND VPWR VPWR _20808_/Y sky130_fd_sc_hd__nor2_4
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12580_/X _12583_/X _12586_/X _12590_/D VGND VGND VPWR VPWR _12590_/X sky130_fd_sc_hd__or4_4
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24576_ _25084_/CLK _24576_/D HRESETn VGND VGND VPWR VPWR _24576_/Q sky130_fd_sc_hd__dfrtp_4
X_21788_ _21777_/A _19515_/Y _14529_/X VGND VGND VPWR VPWR _21788_/X sky130_fd_sc_hd__o21a_4
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20125__A3 _18000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _11518_/Y VGND VGND VPWR VPWR _11541_/X sky130_fd_sc_hd__buf_2
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23527_ _23537_/CLK _23527_/D VGND VGND VPWR VPWR _18895_/A sky130_fd_sc_hd__dfxtp_4
X_20739_ _20739_/A _20739_/B VGND VGND VPWR VPWR _20739_/X sky130_fd_sc_hd__and2_4
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ _14248_/Y VGND VGND VPWR VPWR _14260_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23458_ _24733_/CLK _23458_/D VGND VGND VPWR VPWR _23458_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13211_ _13090_/X _13209_/X _13210_/X VGND VGND VPWR VPWR _13211_/X sky130_fd_sc_hd__and3_4
XFILLER_52_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22409_ _16522_/Y _22488_/B VGND VGND VPWR VPWR _22409_/X sky130_fd_sc_hd__and2_4
X_14191_ _14174_/Y _14190_/X _11980_/A _14150_/X VGND VGND VPWR VPWR _24825_/D sky130_fd_sc_hd__o22a_4
XFILLER_136_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14760__B2 _24107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23389_ _23293_/CLK _23389_/D VGND VGND VPWR VPWR _23389_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_100_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13142_ _13278_/A _13142_/B _13142_/C VGND VGND VPWR VPWR _13142_/X sky130_fd_sc_hd__and3_4
XFILLER_87_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25128_ _25130_/CLK _12215_/Y HRESETn VGND VGND VPWR VPWR _12086_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17973__B _11720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13073_ _13073_/A _13073_/B _13073_/C VGND VGND VPWR VPWR _13073_/X sky130_fd_sc_hd__or3_4
X_17950_ _17918_/A _17948_/X _17950_/C VGND VGND VPWR VPWR _17954_/B sky130_fd_sc_hd__and3_4
XANTENNA__14512__B2 _14484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25059_ _25046_/CLK _25059_/D HRESETn VGND VGND VPWR VPWR _25059_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12024_ _12004_/A _12013_/A _12004_/A _12013_/A VGND VGND VPWR VPWR _12024_/X sky130_fd_sc_hd__a2bb2o_4
X_16901_ _16890_/A _16895_/X _16901_/C VGND VGND VPWR VPWR _16901_/X sky130_fd_sc_hd__and3_4
X_17881_ _17881_/A _23145_/Q VGND VGND VPWR VPWR _17882_/C sky130_fd_sc_hd__or2_4
XFILLER_65_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19620_ _20966_/B _19613_/X _19256_/X _19613_/A VGND VGND VPWR VPWR _23271_/D sky130_fd_sc_hd__a2bb2o_4
X_16832_ _24062_/Q VGND VGND VPWR VPWR _16832_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14276__B1 _14209_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24296__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19551_ _19550_/Y _19546_/X _19256_/X _19533_/Y VGND VGND VPWR VPWR _23295_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16763_ _15908_/Y _24059_/Q _15908_/Y _24059_/Q VGND VGND VPWR VPWR _16764_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13975_ _13974_/X VGND VGND VPWR VPWR _13975_/Y sky130_fd_sc_hd__inv_2
X_18502_ _18502_/A VGND VGND VPWR VPWR _18503_/B sky130_fd_sc_hd__inv_2
XANTENNA__17214__B1 _16671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24225__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15714_ _24466_/Q VGND VGND VPWR VPWR _15717_/C sky130_fd_sc_hd__inv_2
X_12926_ _12925_/X VGND VGND VPWR VPWR _12952_/A sky130_fd_sc_hd__buf_2
X_19482_ _13284_/B VGND VGND VPWR VPWR _19482_/Y sky130_fd_sc_hd__inv_2
X_16694_ _22706_/A _16692_/Y _24387_/Q _17515_/D VGND VGND VPWR VPWR _16694_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18962__B1 _18938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18433_ _23829_/Q VGND VGND VPWR VPWR _18434_/D sky130_fd_sc_hd__inv_2
XFILLER_33_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15645_ _15459_/A _16127_/A VGND VGND VPWR VPWR _15645_/X sky130_fd_sc_hd__or2_4
XANTENNA__15776__B1 _15775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12857_ _25008_/Q VGND VGND VPWR VPWR _12858_/A sky130_fd_sc_hd__inv_2
XANTENNA__12638__A _24462_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21849__B1 _25195_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11808_ _11809_/B _11804_/Y _11815_/C _11804_/Y VGND VGND VPWR VPWR _25181_/D sky130_fd_sc_hd__a2bb2o_4
X_18364_ _16413_/A _23837_/Q _16413_/Y _18363_/Y VGND VGND VPWR VPWR _18364_/X sky130_fd_sc_hd__o22a_4
X_12788_ _22854_/A VGND VGND VPWR VPWR _12788_/Y sky130_fd_sc_hd__inv_2
X_15576_ _15575_/X VGND VGND VPWR VPWR _15576_/X sky130_fd_sc_hd__buf_2
XFILLER_72_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17315_/A VGND VGND VPWR VPWR _17315_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22773__C _22773_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11739_ _11733_/X _11738_/A _11737_/Y _11738_/Y VGND VGND VPWR VPWR _11745_/A sky130_fd_sc_hd__o22a_4
X_14527_ _14448_/B _14526_/Y _14524_/D _14526_/Y VGND VGND VPWR VPWR _14527_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18295_ _18295_/A _18295_/B VGND VGND VPWR VPWR _18296_/C sky130_fd_sc_hd__or2_4
XANTENNA__22827__A1_N _12451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17246_ _17246_/A VGND VGND VPWR VPWR _17246_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23860__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14458_ _14548_/A VGND VGND VPWR VPWR _14544_/A sky130_fd_sc_hd__inv_2
XANTENNA__25084__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19809__A3 _19808_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13409_ _24934_/Q VGND VGND VPWR VPWR _22214_/A sky130_fd_sc_hd__inv_2
XFILLER_31_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14389_ _14368_/Y _14371_/X _14387_/X _24768_/Q _14388_/Y VGND VGND VPWR VPWR _14389_/X
+ sky130_fd_sc_hd__a32o_4
X_17177_ _20372_/A _17176_/X VGND VGND VPWR VPWR _20374_/A sky130_fd_sc_hd__or2_4
XFILLER_116_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25013__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16128_ _15641_/X _16135_/B _15912_/X _20736_/A _16127_/X VGND VGND VPWR VPWR _16128_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22026__B1 _20331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15684__A _15657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16059_ _16071_/A VGND VGND VPWR VPWR _16059_/X sky130_fd_sc_hd__buf_2
XANTENNA__15700__B1 _15386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14503__B2 _14484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22577__A1 _24273_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20588__B1 _20583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19818_ _19818_/A VGND VGND VPWR VPWR _19818_/X sky130_fd_sc_hd__buf_2
XFILLER_110_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19749_ _19749_/A VGND VGND VPWR VPWR _21349_/B sky130_fd_sc_hd__inv_2
XFILLER_65_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22310__A _14047_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22760_ _24452_/Q _22703_/B VGND VGND VPWR VPWR _22760_/X sky130_fd_sc_hd__or2_4
XFILLER_37_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21552__A2 _16134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21711_ _15322_/A _21710_/X _21058_/X _24400_/Q _22148_/A VGND VGND VPWR VPWR _21712_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_80_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22691_ _22691_/A _22688_/X _22691_/C VGND VGND VPWR VPWR _22718_/A sky130_fd_sc_hd__and3_4
XFILLER_129_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22964__B _22959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24430_ _24372_/CLK _15803_/X HRESETn VGND VGND VPWR VPWR _21055_/A sky130_fd_sc_hd__dfrtp_4
X_21642_ _20800_/X VGND VGND VPWR VPWR _21642_/X sky130_fd_sc_hd__buf_2
XANTENNA__23948__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21304__A2 _13357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15782__A3 _16087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15519__B1 _15393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15859__A _24414_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24361_ _24361_/CLK _24361_/D HRESETn VGND VGND VPWR VPWR _21044_/A sky130_fd_sc_hd__dfrtp_4
X_21573_ _24259_/Q _21860_/B VGND VGND VPWR VPWR _21573_/X sky130_fd_sc_hd__and2_4
X_23312_ _23135_/CLK _23312_/D VGND VGND VPWR VPWR _23312_/Q sky130_fd_sc_hd__dfxtp_4
X_20524_ _20524_/A _20524_/B VGND VGND VPWR VPWR _20524_/Y sky130_fd_sc_hd__nor2_4
XFILLER_21_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16192__B1 _16100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24292_ _24590_/CLK _16212_/X HRESETn VGND VGND VPWR VPWR _24292_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23243_ _23258_/CLK _19697_/X VGND VGND VPWR VPWR _19696_/A sky130_fd_sc_hd__dfxtp_4
X_20455_ _15383_/Y _20437_/X _20446_/X _20454_/Y VGND VGND VPWR VPWR _20456_/A sky130_fd_sc_hd__o22a_4
XFILLER_88_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23174_ _23332_/CLK _23174_/D VGND VGND VPWR VPWR _19882_/A sky130_fd_sc_hd__dfxtp_4
X_20386_ _20389_/B _20386_/B _20373_/X VGND VGND VPWR VPWR _20386_/X sky130_fd_sc_hd__and3_4
XFILLER_137_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22125_ _22677_/A _22124_/X VGND VGND VPWR VPWR _22125_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_102_0_HCLK clkbuf_7_51_0_HCLK/X VGND VGND VPWR VPWR _24618_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_133_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22568__B2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24736__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_165_0_HCLK clkbuf_7_82_0_HCLK/X VGND VGND VPWR VPWR _25050_/CLK sky130_fd_sc_hd__clkbuf_1
X_22056_ _22055_/X _22056_/B VGND VGND VPWR VPWR _22056_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_8_0_HCLK clkbuf_6_4_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21007_ _21007_/A _21005_/X _21006_/X VGND VGND VPWR VPWR _21007_/X sky130_fd_sc_hd__and3_4
XFILLER_88_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17444__B1 _17345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14258__B1 _14221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19197__B1 _19152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13760_ _13753_/C VGND VGND VPWR VPWR _13761_/A sky130_fd_sc_hd__buf_2
X_22958_ _24574_/Q _22557_/X _22558_/X _22957_/X VGND VGND VPWR VPWR _22958_/X sky130_fd_sc_hd__a211o_4
XFILLER_21_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16353__A1_N _16351_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22740__B2 _22170_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12711_ _12565_/Y _12716_/B _12666_/X VGND VGND VPWR VPWR _12711_/Y sky130_fd_sc_hd__a21oi_4
X_21909_ _21924_/A _21909_/B VGND VGND VPWR VPWR _21909_/X sky130_fd_sc_hd__or2_4
XFILLER_44_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13691_ _13678_/X _13691_/B VGND VGND VPWR VPWR _13691_/X sky130_fd_sc_hd__or2_4
XANTENNA__15758__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22889_ _22195_/X _22888_/X _22629_/X _12089_/A _22198_/X VGND VGND VPWR VPWR _22890_/B
+ sky130_fd_sc_hd__a32o_4
X_12642_ _12605_/Y _12612_/Y VGND VGND VPWR VPWR _12642_/X sky130_fd_sc_hd__or2_4
X_15430_ _15430_/A VGND VGND VPWR VPWR _15430_/X sky130_fd_sc_hd__buf_2
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23689__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24628_ _23676_/CLK _15283_/X HRESETn VGND VGND VPWR VPWR _24628_/Q sky130_fd_sc_hd__dfstp_4
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15361_ _15361_/A VGND VGND VPWR VPWR _15361_/Y sky130_fd_sc_hd__inv_2
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ _25061_/Q _24526_/Q _12571_/Y _12572_/Y VGND VGND VPWR VPWR _12577_/C sky130_fd_sc_hd__o22a_4
XANTENNA__23618__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24559_ _24545_/CLK _15500_/X HRESETn VGND VGND VPWR VPWR _24559_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21846__A3 _21432_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17100_ _16968_/Y _17097_/X VGND VGND VPWR VPWR _17100_/X sky130_fd_sc_hd__or2_4
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11524_ _25219_/Q VGND VGND VPWR VPWR _11524_/Y sky130_fd_sc_hd__inv_2
X_14312_ _14311_/X VGND VGND VPWR VPWR _14312_/Y sky130_fd_sc_hd__inv_2
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15292_ _15290_/Y _15285_/X _15291_/X _15285_/A VGND VGND VPWR VPWR _15292_/X sky130_fd_sc_hd__a2bb2o_4
X_18080_ _18080_/A VGND VGND VPWR VPWR _18080_/Y sky130_fd_sc_hd__inv_2
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22890__A _22681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14243_ _14226_/A VGND VGND VPWR VPWR _14243_/X sky130_fd_sc_hd__buf_2
X_17031_ _17031_/A VGND VGND VPWR VPWR _17032_/D sky130_fd_sc_hd__inv_2
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15930__B1 _15753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12744__B1 _12666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14174_ _14150_/X VGND VGND VPWR VPWR _14174_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_61_0_HCLK clkbuf_7_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_61_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_13125_ _13065_/X _13125_/B _13125_/C VGND VGND VPWR VPWR _13125_/X sky130_fd_sc_hd__and3_4
XFILLER_124_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18982_ _18982_/A VGND VGND VPWR VPWR _18982_/X sky130_fd_sc_hd__buf_2
XANTENNA__12921__A _12921_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22114__B _20940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24477__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13056_ _13036_/X _13052_/X _13054_/X _25003_/Q _13057_/A VGND VGND VPWR VPWR _13056_/X
+ sky130_fd_sc_hd__a32o_4
X_17933_ _17716_/X _17931_/X _17933_/C VGND VGND VPWR VPWR _17937_/B sky130_fd_sc_hd__and3_4
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12007_ _11990_/A VGND VGND VPWR VPWR _12007_/X sky130_fd_sc_hd__buf_2
XANTENNA__24406__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17864_ _17928_/A _17864_/B VGND VGND VPWR VPWR _17864_/X sky130_fd_sc_hd__or2_4
XFILLER_94_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19603_ _19603_/A VGND VGND VPWR VPWR _19603_/X sky130_fd_sc_hd__buf_2
X_16815_ _16940_/A VGND VGND VPWR VPWR _16867_/A sky130_fd_sc_hd__buf_2
X_17795_ _17927_/A _18882_/A VGND VGND VPWR VPWR _17795_/X sky130_fd_sc_hd__or2_4
XANTENNA__22130__A _24474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19534_ _19533_/Y VGND VGND VPWR VPWR _19534_/X sky130_fd_sc_hd__buf_2
XANTENNA__17224__A _11728_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16746_ _16746_/A _16745_/X VGND VGND VPWR VPWR _16746_/X sky130_fd_sc_hd__or2_4
X_13958_ _13952_/X _13957_/X _13924_/A _13952_/X VGND VGND VPWR VPWR _24894_/D sky130_fd_sc_hd__a2bb2o_4
X_12909_ _12779_/Y _12907_/A VGND VGND VPWR VPWR _12910_/C sky130_fd_sc_hd__or2_4
X_19465_ _20993_/B _19458_/X _18662_/X _19440_/Y VGND VGND VPWR VPWR _19465_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15749__B1 _24459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16677_ _14563_/A VGND VGND VPWR VPWR _17725_/A sky130_fd_sc_hd__inv_2
X_13889_ _20164_/A VGND VGND VPWR VPWR _13890_/A sky130_fd_sc_hd__inv_2
X_18416_ _18472_/A VGND VGND VPWR VPWR _18416_/Y sky130_fd_sc_hd__inv_2
X_15628_ _15604_/A VGND VGND VPWR VPWR _15628_/X sky130_fd_sc_hd__buf_2
X_19396_ _19396_/A VGND VGND VPWR VPWR _19396_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15764__A3 _15600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18347_ _18347_/A _18347_/B _18344_/X _18347_/D VGND VGND VPWR VPWR _18347_/X sky130_fd_sc_hd__or4_4
XFILLER_33_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15559_ _19455_/A VGND VGND VPWR VPWR _15559_/X sky130_fd_sc_hd__buf_2
X_18278_ _18278_/A _18277_/X VGND VGND VPWR VPWR _18282_/B sky130_fd_sc_hd__or2_4
XANTENNA__23039__A2 _21651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16713__A2 _22202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17229_ _11738_/A _17228_/A _11738_/Y _17228_/Y VGND VGND VPWR VPWR _17233_/C sky130_fd_sc_hd__o22a_4
XANTENNA__22247__B1 _24405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11538__A1 _11533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22798__A1 _15572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19112__B1 _19089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20240_ _20244_/A _20239_/X _20212_/B VGND VGND VPWR VPWR _20240_/X sky130_fd_sc_hd__o21a_4
XFILLER_131_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20171_ _23779_/Q _20171_/B VGND VGND VPWR VPWR _20196_/A sky130_fd_sc_hd__and2_4
XFILLER_115_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15515__A1_N _12098_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22024__B _22024_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_238_0_HCLK clkbuf_8_239_0_HCLK/A VGND VGND VPWR VPWR _23753_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24147__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23930_ _24735_/CLK _23930_/D HRESETn VGND VGND VPWR VPWR _23930_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22970__A1 _22335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22970__B2 _22840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23861_ _23762_/CLK _18284_/X HRESETn VGND VGND VPWR VPWR _23861_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15988__B1 _15894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20981__B1 _20968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22812_ _22811_/X VGND VGND VPWR VPWR _22812_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23792_ _24840_/CLK _14151_/Y HRESETn VGND VGND VPWR VPWR _12053_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_38_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22743_ _22734_/X _22743_/B _22743_/C VGND VGND VPWR VPWR _22743_/X sky130_fd_sc_hd__or3_4
XFILLER_0_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23782__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22674_ _24047_/Q _22956_/B VGND VGND VPWR VPWR _22674_/X sky130_fd_sc_hd__or2_4
XFILLER_16_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24413_ _24412_/CLK _24413_/D HRESETn VGND VGND VPWR VPWR _15862_/A sky130_fd_sc_hd__dfrtp_4
X_21625_ _21625_/A _19654_/Y VGND VGND VPWR VPWR _21625_/X sky130_fd_sc_hd__or2_4
XANTENNA__23711__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24344_ _24225_/CLK _16074_/X HRESETn VGND VGND VPWR VPWR _24344_/Q sky130_fd_sc_hd__dfrtp_4
X_21556_ _20221_/B _14016_/X _14055_/A _20744_/X VGND VGND VPWR VPWR _21556_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20507_ _20513_/B VGND VGND VPWR VPWR _20508_/A sky130_fd_sc_hd__inv_2
XANTENNA__24988__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24275_ _24681_/CLK _16260_/X HRESETn VGND VGND VPWR VPWR _24275_/Q sky130_fd_sc_hd__dfrtp_4
X_21487_ _21483_/X _21486_/X _21172_/X VGND VGND VPWR VPWR _21487_/X sky130_fd_sc_hd__o21a_4
XFILLER_106_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22789__B2 _21576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24917__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23226_ _23112_/CLK _19748_/X VGND VGND VPWR VPWR _19747_/A sky130_fd_sc_hd__dfxtp_4
X_20438_ _20438_/A VGND VGND VPWR VPWR _20438_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22215__A _22215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_48_0_HCLK clkbuf_6_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_48_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23157_ _23154_/CLK _23157_/D VGND VGND VPWR VPWR _19929_/A sky130_fd_sc_hd__dfxtp_4
X_20369_ _17176_/X _20369_/B _20349_/X VGND VGND VPWR VPWR _20369_/X sky130_fd_sc_hd__and3_4
XFILLER_79_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22108_ _20967_/A _22108_/B _22107_/X VGND VGND VPWR VPWR _22108_/X sky130_fd_sc_hd__and3_4
XANTENNA__24570__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23088_ _23288_/CLK _23088_/D VGND VGND VPWR VPWR _23088_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_103_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22869__B _22933_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14930_ _24668_/Q _24273_/Q _15106_/A _14929_/Y VGND VGND VPWR VPWR _14931_/D sky130_fd_sc_hd__o22a_4
X_22039_ _22034_/X _22039_/B _22037_/X _22038_/X VGND VGND VPWR VPWR _22039_/X sky130_fd_sc_hd__or4_4
XFILLER_88_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13365__A1_N _11904_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22961__B2 _22322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14861_ _24708_/Q _14859_/Y _24702_/Q _14860_/Y VGND VGND VPWR VPWR _14862_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16600_ _16581_/X _16597_/X _16096_/A _24137_/Q _16590_/X VGND VGND VPWR VPWR _16600_/X
+ sky130_fd_sc_hd__a32o_4
X_13812_ _24899_/Q _24898_/Q VGND VGND VPWR VPWR _13812_/X sky130_fd_sc_hd__or2_4
XANTENNA__17044__A _17124_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_3_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_6_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17580_ _22395_/A _17580_/B VGND VGND VPWR VPWR _17580_/X sky130_fd_sc_hd__or2_4
XFILLER_63_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14792_ _15078_/A _24099_/Q _14791_/X _24096_/Q VGND VGND VPWR VPWR _14792_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16531_ _22282_/A _16530_/X _16279_/X _16530_/X VGND VGND VPWR VPWR _16531_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13743_ _13743_/A VGND VGND VPWR VPWR _14074_/A sky130_fd_sc_hd__inv_2
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19250_ _19250_/A VGND VGND VPWR VPWR _19250_/Y sky130_fd_sc_hd__inv_2
X_16462_ _16462_/A VGND VGND VPWR VPWR _16462_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13674_ _13421_/Y _13671_/X _13398_/X _13671_/X VGND VGND VPWR VPWR _24926_/D sky130_fd_sc_hd__a2bb2o_4
X_18201_ _18200_/Y _18240_/C VGND VGND VPWR VPWR _18201_/X sky130_fd_sc_hd__or2_4
X_15413_ _15413_/A VGND VGND VPWR VPWR _21280_/A sky130_fd_sc_hd__buf_2
X_12625_ _25067_/Q VGND VGND VPWR VPWR _12657_/A sky130_fd_sc_hd__inv_2
X_19181_ _19181_/A VGND VGND VPWR VPWR _19181_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15499__A _11585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16393_ _16043_/A _23763_/Q _16041_/X _16393_/D VGND VGND VPWR VPWR _16393_/X sky130_fd_sc_hd__and4_4
XANTENNA__14954__B2 _14897_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11768__A1 _21188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19342__B1 _19227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18132_ _16098_/Y _18212_/A _16098_/Y _18212_/A VGND VGND VPWR VPWR _18132_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12556_ _24512_/Q VGND VGND VPWR VPWR _12556_/Y sky130_fd_sc_hd__inv_2
X_15344_ _24607_/Q VGND VGND VPWR VPWR _22753_/A sky130_fd_sc_hd__inv_2
XANTENNA__16156__B1 _15479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11507_ _11507_/A _20842_/B VGND VGND VPWR VPWR _11507_/X sky130_fd_sc_hd__or2_4
X_18063_ _11734_/Y VGND VGND VPWR VPWR _18968_/A sky130_fd_sc_hd__buf_2
XFILLER_89_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12487_ _12489_/B VGND VGND VPWR VPWR _12487_/Y sky130_fd_sc_hd__inv_2
X_15275_ _20393_/A VGND VGND VPWR VPWR _15275_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15903__B1 _15282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17014_ _16140_/Y _17021_/A _16140_/Y _17021_/A VGND VGND VPWR VPWR _17017_/B sky130_fd_sc_hd__a2bb2o_4
X_14226_ _14226_/A VGND VGND VPWR VPWR _14226_/X sky130_fd_sc_hd__buf_2
XANTENNA__24658__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22125__A _22677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14157_ _12048_/A VGND VGND VPWR VPWR _14160_/A sky130_fd_sc_hd__inv_2
XFILLER_98_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13108_ _11743_/A _23341_/Q VGND VGND VPWR VPWR _13108_/X sky130_fd_sc_hd__or2_4
X_14088_ _24858_/Q VGND VGND VPWR VPWR _14088_/Y sky130_fd_sc_hd__inv_2
X_18965_ _18963_/Y _18958_/X _18964_/X _18958_/A VGND VGND VPWR VPWR _18965_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22779__B _22147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24240__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13039_ _13042_/A _13039_/B VGND VGND VPWR VPWR _13040_/C sky130_fd_sc_hd__or2_4
X_17916_ _17916_/A _23432_/Q VGND VGND VPWR VPWR _17918_/B sky130_fd_sc_hd__or2_4
XFILLER_26_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18896_ _18895_/Y _18891_/X _18828_/X _18876_/Y VGND VGND VPWR VPWR _23527_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17847_ _17879_/A _17845_/X _17846_/X VGND VGND VPWR VPWR _17851_/B sky130_fd_sc_hd__and3_4
XFILLER_94_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14578__A _14577_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_68_0_HCLK clkbuf_8_69_0_HCLK/A VGND VGND VPWR VPWR _23796_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15434__A2 _15415_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17778_ _17816_/A _23436_/Q VGND VGND VPWR VPWR _17778_/X sky130_fd_sc_hd__or2_4
XFILLER_19_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19517_ _19515_/Y _19511_/X _19448_/X _19516_/X VGND VGND VPWR VPWR _19517_/X sky130_fd_sc_hd__a2bb2o_4
X_16729_ _15957_/Y _16718_/A _22706_/A _16692_/Y VGND VGND VPWR VPWR _16729_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11714__B _11711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24968__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19448_ _19448_/A VGND VGND VPWR VPWR _19448_/X sky130_fd_sc_hd__buf_2
XANTENNA__15737__A3 _15735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21204__A _21374_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19379_ _19377_/Y _19373_/X _19311_/X _19378_/X VGND VGND VPWR VPWR _23356_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14945__B2 _22399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21410_ _20815_/X _21410_/B VGND VGND VPWR VPWR _21410_/X sky130_fd_sc_hd__and2_4
X_22390_ _22390_/A VGND VGND VPWR VPWR _22390_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16698__A1 _22598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21341_ _20965_/A VGND VGND VPWR VPWR _21342_/A sky130_fd_sc_hd__buf_2
XANTENNA__21858__B _21720_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24399__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24060_ _24618_/CLK _24060_/D HRESETn VGND VGND VPWR VPWR _24060_/Q sky130_fd_sc_hd__dfrtp_4
X_21272_ _21265_/X _21271_/X _21062_/X VGND VGND VPWR VPWR _21272_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15370__A1 _15368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23011_ _22919_/A _23001_/X _23004_/X _23010_/X VGND VGND VPWR VPWR _23011_/X sky130_fd_sc_hd__or4_4
X_20223_ _20222_/X VGND VGND VPWR VPWR _20266_/C sky130_fd_sc_hd__inv_2
XANTENNA__24328__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17129__A _17129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20154_ _15297_/X VGND VGND VPWR VPWR _20155_/B sky130_fd_sc_hd__inv_2
XFILLER_98_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15872__A _24409_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20085_ _20084_/Y _20082_/X _19607_/A _20082_/X VGND VGND VPWR VPWR _23098_/D sky130_fd_sc_hd__a2bb2o_4
X_24962_ _24962_/CLK _13570_/X HRESETn VGND VGND VPWR VPWR _13549_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20549__A3 _13515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23913_ _24928_/CLK _18001_/X HRESETn VGND VGND VPWR VPWR _23913_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18396__A1_N _16464_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24893_ _24783_/CLK _24893_/D HRESETn VGND VGND VPWR VPWR _13939_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13436__A1 _24932_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23963__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23844_ _23824_/CLK _23844_/D HRESETn VGND VGND VPWR VPWR _23844_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25187__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17799__A _14571_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23775_ _24897_/CLK _23775_/D HRESETn VGND VGND VPWR VPWR _20163_/C sky130_fd_sc_hd__dfrtp_4
X_20987_ _22105_/A _20986_/X _23941_/Q VGND VGND VPWR VPWR _20987_/X sky130_fd_sc_hd__a21o_4
XANTENNA__25116__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20937__B _20900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16386__B1 _16216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22726_ _22725_/X VGND VGND VPWR VPWR _22744_/B sky130_fd_sc_hd__inv_2
XFILLER_129_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22657_ _21069_/X VGND VGND VPWR VPWR _22657_/X sky130_fd_sc_hd__buf_2
XANTENNA__19324__B1 _19232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12410_ _12469_/A VGND VGND VPWR VPWR _12410_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11640__A _25190_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21608_ _21612_/A _21608_/B VGND VGND VPWR VPWR _21610_/B sky130_fd_sc_hd__or2_4
XFILLER_51_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13390_ _14106_/B VGND VGND VPWR VPWR _13390_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_11_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22588_ _22011_/X _22586_/X _22322_/X _22587_/X VGND VGND VPWR VPWR _22588_/X sky130_fd_sc_hd__o22a_4
X_12341_ _12432_/A VGND VGND VPWR VPWR _12433_/A sky130_fd_sc_hd__inv_2
X_21539_ _20837_/X VGND VGND VPWR VPWR _22943_/A sky130_fd_sc_hd__buf_2
XANTENNA__16689__B2 _17498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24327_ _23852_/CLK _16120_/X HRESETn VGND VGND VPWR VPWR _24327_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15060_ _14869_/B _15059_/X VGND VGND VPWR VPWR _15061_/B sky130_fd_sc_hd__or2_4
XANTENNA__24751__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12272_ _12275_/A _12278_/B VGND VGND VPWR VPWR _12276_/B sky130_fd_sc_hd__or2_4
XFILLER_107_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24258_ _24259_/CLK _16289_/X HRESETn VGND VGND VPWR VPWR _24258_/Q sky130_fd_sc_hd__dfrtp_4
X_14011_ _14010_/X VGND VGND VPWR VPWR _24880_/D sky130_fd_sc_hd__inv_2
XANTENNA__24069__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23209_ _23303_/CLK _19794_/X VGND VGND VPWR VPWR _19792_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24024__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24189_ _24167_/CLK _24189_/D HRESETn VGND VGND VPWR VPWR _24189_/Q sky130_fd_sc_hd__dfrtp_4
X_18750_ _18749_/Y _18745_/X _18679_/X _18745_/X VGND VGND VPWR VPWR _23578_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16689__A2_N _17498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15962_ _15959_/Y _15961_/X _11576_/X _15961_/X VGND VGND VPWR VPWR _15962_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_221_0_HCLK clkbuf_8_221_0_HCLK/A VGND VGND VPWR VPWR _23830_/CLK sky130_fd_sc_hd__clkbuf_1
X_17701_ _17698_/A _17701_/B VGND VGND VPWR VPWR _17701_/X sky130_fd_sc_hd__or2_4
XFILLER_88_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14913_ _24279_/Q VGND VGND VPWR VPWR _14913_/Y sky130_fd_sc_hd__inv_2
X_18681_ _23601_/Q VGND VGND VPWR VPWR _18681_/Y sky130_fd_sc_hd__inv_2
X_15893_ _15885_/A VGND VGND VPWR VPWR _15893_/X sky130_fd_sc_hd__buf_2
XFILLER_114_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17632_ _17632_/A VGND VGND VPWR VPWR _17632_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14844_ _14844_/A VGND VGND VPWR VPWR _15067_/C sky130_fd_sc_hd__buf_2
XFILLER_90_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17563_ _16697_/Y _17563_/B VGND VGND VPWR VPWR _17563_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__23633__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14775_ _14809_/A _24115_/Q _24692_/Q _14709_/Y VGND VGND VPWR VPWR _14784_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11987_ _11986_/X VGND VGND VPWR VPWR _21564_/A sky130_fd_sc_hd__buf_2
X_19302_ _13023_/B VGND VGND VPWR VPWR _19302_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16514_ _16513_/Y _16511_/X _16266_/X _16511_/X VGND VGND VPWR VPWR _24175_/D sky130_fd_sc_hd__a2bb2o_4
X_13726_ _24640_/Q VGND VGND VPWR VPWR _13726_/X sky130_fd_sc_hd__buf_2
X_17494_ _22376_/A VGND VGND VPWR VPWR _17494_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16377__B1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19233_ _19231_/Y _19226_/X _19232_/X _19212_/Y VGND VGND VPWR VPWR _23407_/D sky130_fd_sc_hd__a2bb2o_4
X_16445_ _24201_/Q VGND VGND VPWR VPWR _16445_/Y sky130_fd_sc_hd__inv_2
X_13657_ _13649_/A VGND VGND VPWR VPWR _13657_/X sky130_fd_sc_hd__buf_2
XFILLER_31_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19315__B1 _19221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11550__A _25214_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12608_ _12607_/Y _24519_/Q _25058_/Q _12559_/Y VGND VGND VPWR VPWR _12608_/X sky130_fd_sc_hd__a2bb2o_4
X_19164_ _17948_/B VGND VGND VPWR VPWR _19164_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24839__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16376_ _16376_/A VGND VGND VPWR VPWR _16376_/X sky130_fd_sc_hd__buf_2
XFILLER_121_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13588_ _13562_/X _13580_/X _13585_/Y _13587_/X _11685_/A VGND VGND VPWR VPWR _13588_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20863__A _20863_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18115_ _18115_/A VGND VGND VPWR VPWR _21898_/A sky130_fd_sc_hd__inv_2
X_15327_ _15353_/A VGND VGND VPWR VPWR _15327_/X sky130_fd_sc_hd__buf_2
X_12539_ _12456_/X _12536_/B _12539_/C VGND VGND VPWR VPWR _12539_/X sky130_fd_sc_hd__and3_4
X_19095_ _18801_/X VGND VGND VPWR VPWR _19095_/X sky130_fd_sc_hd__buf_2
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24492__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18046_ _21335_/A _18022_/X _21335_/A _18022_/X VGND VGND VPWR VPWR _18046_/X sky130_fd_sc_hd__a2bb2o_4
X_15258_ _14100_/X _23764_/Q _15251_/Y _13716_/C _15254_/X VGND VGND VPWR VPWR _15258_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_32_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24421__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14209_ _13632_/A VGND VGND VPWR VPWR _14209_/X sky130_fd_sc_hd__buf_2
XFILLER_98_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15189_ _15191_/B VGND VGND VPWR VPWR _15190_/B sky130_fd_sc_hd__inv_2
XFILLER_28_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21694__A _22870_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_31_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19997_ _19995_/Y _19991_/X _19424_/X _19996_/X VGND VGND VPWR VPWR _23132_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18948_ _18947_/Y _18945_/X _18880_/X _18945_/X VGND VGND VPWR VPWR _18948_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21189__B1 _20745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18879_ _23533_/Q VGND VGND VPWR VPWR _18879_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20910_ _20909_/X VGND VGND VPWR VPWR _20910_/X sky130_fd_sc_hd__buf_2
X_21890_ _21886_/X _21890_/B VGND VGND VPWR VPWR _21890_/Y sky130_fd_sc_hd__nor2_4
XFILLER_66_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20841_ _17222_/B VGND VGND VPWR VPWR _20842_/C sky130_fd_sc_hd__inv_2
XPHY_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23560_ _23560_/CLK _23560_/D VGND VGND VPWR VPWR _18800_/A sky130_fd_sc_hd__dfxtp_4
X_20772_ _20772_/A VGND VGND VPWR VPWR _20772_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22511_ _22510_/X VGND VGND VPWR VPWR _22997_/A sky130_fd_sc_hd__inv_2
XFILLER_74_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23491_ _23493_/CLK _23491_/D VGND VGND VPWR VPWR _23491_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15040__B1 _15027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19306__B1 _19170_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22972__B _22015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22442_ _16438_/Y _20833_/X _21715_/X _22441_/X VGND VGND VPWR VPWR _22443_/A sky130_fd_sc_hd__a211o_4
XANTENNA__20773__A _11514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24509__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25161_ _23885_/CLK _25161_/D HRESETn VGND VGND VPWR VPWR _11926_/A sky130_fd_sc_hd__dfrtp_4
X_22373_ _22373_/A _22524_/B VGND VGND VPWR VPWR _22373_/X sky130_fd_sc_hd__or2_4
XANTENNA__22861__B1 _22858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21588__B _21582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_113_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_227_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24112_ _24112_/CLK _24112_/D HRESETn VGND VGND VPWR VPWR _14737_/A sky130_fd_sc_hd__dfrtp_4
X_21324_ _21324_/A _21324_/B _21296_/X _21323_/X VGND VGND VPWR VPWR _21324_/X sky130_fd_sc_hd__or4_4
X_25092_ _25097_/CLK _12463_/Y HRESETn VGND VGND VPWR VPWR _25092_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16540__B1 _16373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13354__B1 _11981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24162__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24043_ _24307_/CLK _24043_/D HRESETn VGND VGND VPWR VPWR _17041_/A sky130_fd_sc_hd__dfrtp_4
X_21255_ _21250_/X _21254_/Y _13421_/Y _21250_/X VGND VGND VPWR VPWR _21255_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20206_ _20202_/Y _20203_/Y _13711_/X _20205_/Y VGND VGND VPWR VPWR _20206_/X sky130_fd_sc_hd__a211o_4
XFILLER_2_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21186_ _21109_/B VGND VGND VPWR VPWR _22198_/A sky130_fd_sc_hd__buf_2
XFILLER_133_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20137_ _20133_/Y _20136_/X _17993_/X _20136_/X VGND VGND VPWR VPWR _23076_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22212__B _22497_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14854__B1 _14997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20068_ _20066_/Y _20060_/X _19808_/X _20067_/X VGND VGND VPWR VPWR _20068_/X sky130_fd_sc_hd__a2bb2o_4
X_24945_ _24071_/CLK _13633_/X HRESETn VGND VGND VPWR VPWR _13622_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_86_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11635__A _11635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11910_ _11910_/A VGND VGND VPWR VPWR _11910_/Y sky130_fd_sc_hd__inv_2
X_12890_ _12890_/A _12890_/B VGND VGND VPWR VPWR _12891_/C sky130_fd_sc_hd__or2_4
X_24876_ _24879_/CLK _14035_/X HRESETn VGND VGND VPWR VPWR _20209_/B sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_51_0_HCLK clkbuf_8_51_0_HCLK/A VGND VGND VPWR VPWR _23986_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11841_ _11838_/Y _11831_/X _11839_/X _11840_/X VGND VGND VPWR VPWR _25174_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23827_ _23828_/CLK _18513_/Y HRESETn VGND VGND VPWR VPWR _23827_/Q sky130_fd_sc_hd__dfrtp_4
X_11772_ _25184_/Q _11772_/B _25185_/Q VGND VGND VPWR VPWR _11773_/C sky130_fd_sc_hd__and3_4
X_14560_ _14560_/A VGND VGND VPWR VPWR _14560_/Y sky130_fd_sc_hd__inv_2
X_23758_ _24168_/CLK _20683_/X HRESETn VGND VGND VPWR VPWR _23758_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13511_ _13510_/X VGND VGND VPWR VPWR _20524_/B sky130_fd_sc_hd__buf_2
X_22709_ _24310_/Q _22897_/B VGND VGND VPWR VPWR _22709_/X sky130_fd_sc_hd__or2_4
X_14491_ _14541_/D _14460_/X _14490_/Y VGND VGND VPWR VPWR _14491_/X sky130_fd_sc_hd__o21a_4
XFILLER_110_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15031__B1 _14984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23689_ _23767_/CLK _20407_/X HRESETn VGND VGND VPWR VPWR _23689_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16230_ _20856_/A VGND VGND VPWR VPWR _22017_/A sky130_fd_sc_hd__buf_2
X_13442_ _13442_/A VGND VGND VPWR VPWR _14424_/B sky130_fd_sc_hd__buf_2
XANTENNA__21779__A _21519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24932__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13373_ _11890_/Y _13372_/X _11626_/X _13372_/X VGND VGND VPWR VPWR _13373_/X sky130_fd_sc_hd__a2bb2o_4
X_16161_ _16160_/Y _16158_/X _15484_/X _16158_/X VGND VGND VPWR VPWR _24312_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15777__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_24_0_HCLK_A clkbuf_4_12_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15112_ _15112_/A _15197_/A _15112_/C _14903_/Y VGND VGND VPWR VPWR _15112_/X sky130_fd_sc_hd__or4_4
X_12324_ _12315_/X _12324_/B _12321_/X _12323_/X VGND VGND VPWR VPWR _12352_/B sky130_fd_sc_hd__or4_4
X_16092_ _24337_/Q VGND VGND VPWR VPWR _22401_/A sky130_fd_sc_hd__inv_2
XANTENNA__16531__B1 _16279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13345__B1 _11620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12255_ _12165_/X VGND VGND VPWR VPWR _12261_/A sky130_fd_sc_hd__buf_2
X_15043_ _15043_/A VGND VGND VPWR VPWR _15044_/B sky130_fd_sc_hd__inv_2
X_19920_ _23160_/Q VGND VGND VPWR VPWR _21229_/B sky130_fd_sc_hd__inv_2
XFILLER_119_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19851_ _23186_/Q VGND VGND VPWR VPWR _21509_/B sky130_fd_sc_hd__inv_2
X_12186_ _12154_/Y _12186_/B _12193_/A _12192_/A VGND VGND VPWR VPWR _12189_/B sky130_fd_sc_hd__or4_4
Xclkbuf_5_18_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18802_ _18801_/X VGND VGND VPWR VPWR _18802_/X sky130_fd_sc_hd__buf_2
X_19782_ _19778_/Y _19781_/X _19442_/X _19781_/X VGND VGND VPWR VPWR _23214_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23885__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16994_ _21066_/A VGND VGND VPWR VPWR _17160_/A sky130_fd_sc_hd__inv_2
XANTENNA__16401__A _16401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18733_ _14581_/A _19123_/B VGND VGND VPWR VPWR _18734_/D sky130_fd_sc_hd__or2_4
XFILLER_27_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15945_ _24382_/Q VGND VGND VPWR VPWR _15945_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23814__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25038__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11545__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18664_ _23606_/Q VGND VGND VPWR VPWR _18664_/Y sky130_fd_sc_hd__inv_2
X_15876_ _15875_/Y _15873_/X _11590_/X _15873_/X VGND VGND VPWR VPWR _24408_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17615_ _17615_/A _17615_/B VGND VGND VPWR VPWR _17615_/X sky130_fd_sc_hd__or2_4
X_14827_ _24138_/Q VGND VGND VPWR VPWR _14827_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18595_ _16351_/Y _23827_/Q _16351_/Y _23827_/Q VGND VGND VPWR VPWR _18595_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17546_ _17545_/X VGND VGND VPWR VPWR _23964_/D sky130_fd_sc_hd__inv_2
X_14758_ _14757_/Y _24105_/Q _14757_/Y _24105_/Q VGND VGND VPWR VPWR _14761_/C sky130_fd_sc_hd__a2bb2o_4
X_13709_ _23687_/Q _13708_/X _14096_/A _13682_/Y VGND VGND VPWR VPWR _13709_/X sky130_fd_sc_hd__o22a_4
X_17477_ _17619_/A VGND VGND VPWR VPWR _17509_/A sky130_fd_sc_hd__buf_2
XANTENNA__21894__B2 _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14689_ _14689_/A VGND VGND VPWR VPWR _24716_/D sky130_fd_sc_hd__inv_2
X_19216_ _19215_/Y _19213_/X _19149_/X _19213_/X VGND VGND VPWR VPWR _23413_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16428_ _24208_/Q VGND VGND VPWR VPWR _16428_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21689__A _20782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24673__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16770__B1 _15846_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19147_ _19143_/Y _19146_/X _19059_/X _19146_/X VGND VGND VPWR VPWR _19147_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24602__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16359_ _16364_/A VGND VGND VPWR VPWR _16359_/X sky130_fd_sc_hd__buf_2
XFILLER_8_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19078_ _18734_/D _18874_/X VGND VGND VPWR VPWR _19078_/Y sky130_fd_sc_hd__nor2_4
XFILLER_133_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12139__B2 _24560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18029_ _18022_/A VGND VGND VPWR VPWR _18038_/A sky130_fd_sc_hd__inv_2
XFILLER_114_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13000__A _12818_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21040_ _22637_/A VGND VGND VPWR VPWR _21040_/X sky130_fd_sc_hd__buf_2
XANTENNA__18275__B1 _18228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17407__A _17303_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22991_ _20545_/Y _20926_/X _20679_/Y _21561_/X VGND VGND VPWR VPWR _22991_/X sky130_fd_sc_hd__o22a_4
XFILLER_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24730_ _24728_/CLK _14632_/X HRESETn VGND VGND VPWR VPWR _24730_/Q sky130_fd_sc_hd__dfrtp_4
X_21942_ _21392_/A _21942_/B VGND VGND VPWR VPWR _21944_/B sky130_fd_sc_hd__or2_4
XFILLER_27_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21871__B _20885_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16589__B1 _24144_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12390__A1_N _12389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_38_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_77_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21873_ _21649_/B _21082_/B _15428_/X _21872_/X VGND VGND VPWR VPWR _21873_/X sky130_fd_sc_hd__a211o_4
X_24661_ _24662_/CLK _24661_/D HRESETn VGND VGND VPWR VPWR _24661_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ _20847_/A VGND VGND VPWR VPWR _21097_/B sky130_fd_sc_hd__buf_2
XPHY_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23612_ _23493_/CLK _23612_/D VGND VGND VPWR VPWR _18649_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24592_ _23734_/CLK _24592_/D HRESETn VGND VGND VPWR VPWR _24592_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22983__A _24123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21885__A1 _25144_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20755_ _13614_/X VGND VGND VPWR VPWR _22036_/A sky130_fd_sc_hd__buf_2
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23543_ _25061_/CLK _23543_/D VGND VGND VPWR VPWR _23543_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23474_ _23471_/CLK _23474_/D VGND VGND VPWR VPWR _13212_/B sky130_fd_sc_hd__dfxtp_4
X_20686_ _11881_/A _20686_/B VGND VGND VPWR VPWR _20686_/Y sky130_fd_sc_hd__nor2_4
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_HCLK clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_22425_ _24481_/Q _22147_/A VGND VGND VPWR VPWR _22425_/X sky130_fd_sc_hd__and2_4
XANTENNA__24343__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25213_ _25214_/CLK _25213_/D HRESETn VGND VGND VPWR VPWR _25213_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22356_ _23922_/Q _12065_/A VGND VGND VPWR VPWR _22356_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__21111__B _11529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25144_ _23789_/CLK _11998_/X HRESETn VGND VGND VPWR VPWR _25144_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21307_ _21072_/X VGND VGND VPWR VPWR _21447_/A sky130_fd_sc_hd__inv_2
XANTENNA__20860__A2 _21093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25075_ _25097_/CLK _12526_/X HRESETn VGND VGND VPWR VPWR _25075_/Q sky130_fd_sc_hd__dfrtp_4
X_22287_ _15463_/A VGND VGND VPWR VPWR _22335_/A sky130_fd_sc_hd__buf_2
X_12040_ _12040_/A VGND VGND VPWR VPWR _12040_/Y sky130_fd_sc_hd__inv_2
X_24026_ _23664_/CLK _17189_/X HRESETn VGND VGND VPWR VPWR _24026_/Q sky130_fd_sc_hd__dfstp_4
X_21238_ _21238_/A VGND VGND VPWR VPWR _21392_/A sky130_fd_sc_hd__buf_2
XFILLER_137_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22223__A _22223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20073__B1 _15416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21169_ _21169_/A _21169_/B VGND VGND VPWR VPWR _21171_/B sky130_fd_sc_hd__or2_4
XANTENNA__23038__B _21807_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16221__A _14369_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13991_ _13952_/A _13990_/Y _24884_/Q _13952_/A VGND VGND VPWR VPWR _24884_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25131__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15730_ _15729_/X VGND VGND VPWR VPWR _15730_/X sky130_fd_sc_hd__buf_2
XFILLER_98_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12942_ _12942_/A VGND VGND VPWR VPWR _25025_/D sky130_fd_sc_hd__inv_2
XFILLER_105_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12358__A1_N _21104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24928_ _24928_/CLK _24928_/D HRESETn VGND VGND VPWR VPWR _24928_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23054__A _23041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15661_ _15661_/A VGND VGND VPWR VPWR _15661_/X sky130_fd_sc_hd__buf_2
X_12873_ _25006_/Q VGND VGND VPWR VPWR _12999_/A sky130_fd_sc_hd__inv_2
XFILLER_2_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24859_ _24859_/CLK _24859_/D HRESETn VGND VGND VPWR VPWR _24859_/Q sky130_fd_sc_hd__dfrtp_4
X_17400_ _17325_/B _17399_/X VGND VGND VPWR VPWR _17400_/X sky130_fd_sc_hd__or2_4
X_14612_ _24723_/Q _14612_/B _14612_/C VGND VGND VPWR VPWR _14612_/X sky130_fd_sc_hd__or3_4
XFILLER_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17052__A _17052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11824_ _11824_/A VGND VGND VPWR VPWR _11824_/Y sky130_fd_sc_hd__inv_2
X_18380_ _24207_/Q _18495_/B _16462_/Y _23818_/Q VGND VGND VPWR VPWR _18380_/X sky130_fd_sc_hd__a2bb2o_4
X_15592_ _12615_/Y _15590_/X _15332_/X _15590_/X VGND VGND VPWR VPWR _15592_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22893__A _22163_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17331_/A VGND VGND VPWR VPWR _17331_/Y sky130_fd_sc_hd__inv_2
X_14543_ _14543_/A VGND VGND VPWR VPWR _14543_/X sky130_fd_sc_hd__buf_2
XPHY_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11755_/A VGND VGND VPWR VPWR _11755_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17262_ _23987_/Q VGND VGND VPWR VPWR _17262_/Y sky130_fd_sc_hd__inv_2
XPHY_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14474_ _19862_/A _14473_/X _19862_/A _14473_/X VGND VGND VPWR VPWR _14474_/X sky130_fd_sc_hd__a2bb2o_4
X_11686_ _13585_/A _22215_/A _13585_/A _22215_/A VGND VGND VPWR VPWR _11693_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19001_ _19000_/Y _18996_/X _15559_/X _18996_/X VGND VGND VPWR VPWR _19001_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16213_ _21293_/A VGND VGND VPWR VPWR _16213_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24084__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13425_ _24939_/Q VGND VGND VPWR VPWR _22449_/A sky130_fd_sc_hd__inv_2
XANTENNA__21302__A _21570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17193_ _17171_/X _17185_/X _20723_/B _24022_/Q _17188_/X VGND VGND VPWR VPWR _17193_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_128_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24809__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22117__B _21543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15300__A _23762_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24013__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16144_ _16137_/A VGND VGND VPWR VPWR _16165_/A sky130_fd_sc_hd__buf_2
X_13356_ _13355_/Y _13351_/X _13330_/X _13338_/Y VGND VGND VPWR VPWR _24987_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16504__B1 _16334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12307_ _24473_/Q VGND VGND VPWR VPWR _12307_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16075_ _16075_/A VGND VGND VPWR VPWR _16075_/Y sky130_fd_sc_hd__inv_2
X_13287_ _11735_/Y _13279_/X _13287_/C VGND VGND VPWR VPWR _13287_/X sky130_fd_sc_hd__and3_4
X_15026_ _15018_/X _15024_/X _15026_/C VGND VGND VPWR VPWR _24703_/D sky130_fd_sc_hd__and3_4
X_19903_ _19903_/A VGND VGND VPWR VPWR _22079_/B sky130_fd_sc_hd__inv_2
X_12238_ _12173_/C _12237_/X VGND VGND VPWR VPWR _12252_/B sky130_fd_sc_hd__or2_4
XANTENNA__22133__A _22133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25219__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12169_ _25130_/Q VGND VGND VPWR VPWR _12170_/B sky130_fd_sc_hd__inv_2
X_19834_ _23192_/Q VGND VGND VPWR VPWR _19834_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16131__A _11944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18009__B1 _16546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16977_ _24051_/Q VGND VGND VPWR VPWR _17026_/B sky130_fd_sc_hd__inv_2
X_19765_ _19759_/Y VGND VGND VPWR VPWR _19765_/X sky130_fd_sc_hd__buf_2
XFILLER_81_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15491__B1 _11566_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15928_ _15921_/X VGND VGND VPWR VPWR _15928_/X sky130_fd_sc_hd__buf_2
X_18716_ _23589_/Q VGND VGND VPWR VPWR _18716_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19442__A _19442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19696_ _19696_/A VGND VGND VPWR VPWR _19696_/Y sky130_fd_sc_hd__inv_2
X_18647_ _23613_/Q VGND VGND VPWR VPWR _21949_/B sky130_fd_sc_hd__inv_2
X_15859_ _24414_/Q VGND VGND VPWR VPWR _15859_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24854__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18578_ _24249_/Q _18462_/A _16385_/Y _23814_/Q VGND VGND VPWR VPWR _18581_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17529_ _17503_/B _17511_/B _17503_/A VGND VGND VPWR VPWR _17529_/X sky130_fd_sc_hd__o21a_4
XFILLER_75_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20540_ _20419_/X _20539_/Y _15331_/A _20465_/X VGND VGND VPWR VPWR _23723_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20471_ _20461_/X _20470_/X _24595_/Q _20466_/X VGND VGND VPWR VPWR _20471_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16306__A _16305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22210_ _22584_/A VGND VGND VPWR VPWR _22500_/A sky130_fd_sc_hd__buf_2
XANTENNA__18496__B1 _18449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12142__A2_N _24567_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23190_ _23179_/CLK _23190_/D VGND VGND VPWR VPWR _19839_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_106_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22141_ _11992_/Y _14013_/B _21581_/A VGND VGND VPWR VPWR _22141_/X sky130_fd_sc_hd__o21a_4
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22072_ _21786_/A _22072_/B VGND VGND VPWR VPWR _22073_/C sky130_fd_sc_hd__or2_4
XANTENNA__22044__B2 _21400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14521__A2 _14437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23736__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12532__A1 _12389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21023_ _13624_/Y _21018_/X _13334_/X _21020_/X _21022_/X VGND VGND VPWR VPWR _21024_/A
+ sky130_fd_sc_hd__a2111o_4
XANTENNA__13665__A _13665_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18015__A3 _16558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22974_ _22974_/A VGND VGND VPWR VPWR _22974_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24713_ _24671_/CLK _14981_/X HRESETn VGND VGND VPWR VPWR _24713_/Q sky130_fd_sc_hd__dfrtp_4
X_21925_ _21342_/A _21925_/B VGND VGND VPWR VPWR _21925_/X sky130_fd_sc_hd__or2_4
XFILLER_3_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24595__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24644_ _24644_/CLK _24644_/D HRESETn VGND VGND VPWR VPWR _13716_/A sky130_fd_sc_hd__dfrtp_4
X_21856_ _20940_/X _21838_/Y _21844_/Y _21855_/X VGND VGND VPWR VPWR _21856_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12599__B2 _24514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24524__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _20832_/A VGND VGND VPWR VPWR _20807_/X sky130_fd_sc_hd__buf_2
XFILLER_19_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21787_ _21762_/X _21787_/B VGND VGND VPWR VPWR _21787_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_125_0_HCLK clkbuf_7_62_0_HCLK/X VGND VGND VPWR VPWR _24641_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24575_ _24488_/CLK _15469_/X HRESETn VGND VGND VPWR VPWR _24575_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11540_ HWDATA[27] VGND VGND VPWR VPWR _11540_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_188_0_HCLK clkbuf_7_94_0_HCLK/X VGND VGND VPWR VPWR _24545_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23526_ _23531_/CLK _18902_/X VGND VGND VPWR VPWR _17682_/B sky130_fd_sc_hd__dfxtp_4
X_20738_ _13009_/A _20738_/B VGND VGND VPWR VPWR _20738_/X sky130_fd_sc_hd__and2_4
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22218__A _16042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20669_ _13540_/A _13539_/X _13541_/X VGND VGND VPWR VPWR _20669_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_109_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23457_ _23457_/CLK _23457_/D VGND VGND VPWR VPWR _19091_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_13_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16216__A _16216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ _13137_/A _13210_/B VGND VGND VPWR VPWR _13210_/X sky130_fd_sc_hd__or2_4
X_22408_ _22408_/A _22188_/X VGND VGND VPWR VPWR _22408_/X sky130_fd_sc_hd__and2_4
XANTENNA__22283__A1 _20927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14190_ _24825_/Q _14169_/B _24824_/Q _14165_/B VGND VGND VPWR VPWR _14190_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20961__A _20961_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23388_ _23388_/CLK _23388_/D VGND VGND VPWR VPWR _19288_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_109_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13141_ _13316_/A _13141_/B VGND VGND VPWR VPWR _13142_/C sky130_fd_sc_hd__or2_4
X_25127_ _25084_/CLK _25127_/D HRESETn VGND VGND VPWR VPWR _12078_/A sky130_fd_sc_hd__dfrtp_4
X_22339_ _24267_/Q _22477_/B _22338_/X VGND VGND VPWR VPWR _22339_/X sky130_fd_sc_hd__o21a_4
XFILLER_87_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13072_ _13065_/X _13068_/X _13072_/C VGND VGND VPWR VPWR _13073_/C sky130_fd_sc_hd__and3_4
XFILLER_3_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14512__A2 _14480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22035__B2 _21088_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25058_ _24523_/CLK _25058_/D HRESETn VGND VGND VPWR VPWR _25058_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12023_ _12001_/A _12022_/A _12001_/Y _12022_/Y VGND VGND VPWR VPWR _12023_/X sky130_fd_sc_hd__o22a_4
X_16900_ _16780_/Y _16900_/B VGND VGND VPWR VPWR _16901_/C sky130_fd_sc_hd__nand2_4
XANTENNA__19987__B1 _19859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24009_ _24008_/CLK _24009_/D HRESETn VGND VGND VPWR VPWR _17237_/A sky130_fd_sc_hd__dfrtp_4
X_17880_ _17944_/A _17880_/B VGND VGND VPWR VPWR _17880_/X sky130_fd_sc_hd__or2_4
XFILLER_105_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16831_ _16927_/A _16935_/A _16771_/Y _16831_/D VGND VGND VPWR VPWR _16838_/A sky130_fd_sc_hd__or4_4
XFILLER_66_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15473__B1 _11525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19550_ _23295_/Q VGND VGND VPWR VPWR _19550_/Y sky130_fd_sc_hd__inv_2
X_16762_ _24416_/Q _16760_/Y _24422_/Q _16866_/A VGND VGND VPWR VPWR _16762_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13974_ _13928_/C _13943_/B _13928_/C _13943_/B VGND VGND VPWR VPWR _13974_/X sky130_fd_sc_hd__a2bb2o_4
X_18501_ _18504_/A _18501_/B _18501_/C VGND VGND VPWR VPWR _23831_/D sky130_fd_sc_hd__and3_4
XFILLER_4_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15713_ _15713_/A VGND VGND VPWR VPWR _15713_/X sky130_fd_sc_hd__buf_2
XFILLER_20_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12925_ _12867_/X VGND VGND VPWR VPWR _12925_/X sky130_fd_sc_hd__buf_2
X_19481_ _19479_/Y _19480_/X _19387_/X _19480_/X VGND VGND VPWR VPWR _19481_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16693_ _16693_/A VGND VGND VPWR VPWR _17515_/D sky130_fd_sc_hd__inv_2
XFILLER_98_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18432_ _18430_/Y _18486_/B _18352_/A _18488_/A VGND VGND VPWR VPWR _18432_/X sky130_fd_sc_hd__or4_4
X_15644_ _21795_/B VGND VGND VPWR VPWR _16127_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_21_0_HCLK clkbuf_7_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12856_ _12856_/A _12856_/B _12856_/C _12855_/X VGND VGND VPWR VPWR _12866_/C sky130_fd_sc_hd__or4_4
XFILLER_92_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12850__A1_N _12972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24265__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_84_0_HCLK clkbuf_6_42_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_84_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_11807_ _11807_/A VGND VGND VPWR VPWR _25182_/D sky130_fd_sc_hd__inv_2
X_18363_ _23837_/Q VGND VGND VPWR VPWR _18363_/Y sky130_fd_sc_hd__inv_2
X_15575_ _11949_/Y _24619_/Q _11512_/Y _11514_/A VGND VGND VPWR VPWR _15575_/X sky130_fd_sc_hd__or4_4
XANTENNA__21849__B2 _22198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12787_ _22243_/A VGND VGND VPWR VPWR _12787_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _17246_/Y _17286_/Y _17313_/X VGND VGND VPWR VPWR _17348_/D sky130_fd_sc_hd__or3_4
X_14526_ _14521_/X VGND VGND VPWR VPWR _14526_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15528__A1 _15411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _11738_/A VGND VGND VPWR VPWR _11738_/Y sky130_fd_sc_hd__inv_2
X_18294_ _23858_/Q _18294_/B VGND VGND VPWR VPWR _18296_/B sky130_fd_sc_hd__or2_4
XANTENNA__22773__D _22772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17245_ _25200_/Q _17415_/A _11544_/Y _24004_/Q VGND VGND VPWR VPWR _17245_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21032__A _12356_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14457_ _24740_/Q VGND VGND VPWR VPWR _14548_/A sky130_fd_sc_hd__buf_2
X_11669_ _11669_/A _11664_/X _11666_/X _11668_/X VGND VGND VPWR VPWR _11669_/X sky130_fd_sc_hd__or4_4
XANTENNA__14200__A1 _14199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ _24929_/Q VGND VGND VPWR VPWR _13408_/Y sky130_fd_sc_hd__inv_2
X_17176_ _20368_/A _20368_/B VGND VGND VPWR VPWR _17176_/X sky130_fd_sc_hd__or2_4
XFILLER_116_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14388_ _14387_/X _14369_/X _24946_/Q VGND VGND VPWR VPWR _14388_/Y sky130_fd_sc_hd__o21ai_4
X_16127_ _16127_/A _15822_/X VGND VGND VPWR VPWR _16127_/X sky130_fd_sc_hd__or2_4
XFILLER_127_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13339_ _13338_/Y VGND VGND VPWR VPWR _13339_/X sky130_fd_sc_hd__buf_2
XANTENNA__22981__A1_N _12391_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16058_ _24350_/Q VGND VGND VPWR VPWR _16058_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14503__A2 _14480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22026__B2 _22227_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25053__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15009_ _15014_/A _15009_/B _15008_/X VGND VGND VPWR VPWR _15009_/X sky130_fd_sc_hd__and3_4
XANTENNA__19978__B1 _19452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22577__A2 _22477_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19817_ _19817_/A VGND VGND VPWR VPWR _21957_/B sky130_fd_sc_hd__inv_2
XFILLER_69_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19748_ _21482_/B _19743_/X _19724_/X _19743_/X VGND VGND VPWR VPWR _19748_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21537__B1 _21793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19679_ _23249_/Q VGND VGND VPWR VPWR _19679_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21710_ _24294_/Q _21710_/B VGND VGND VPWR VPWR _21710_/X sky130_fd_sc_hd__or2_4
X_22690_ _24146_/Q _22505_/X _22576_/X _22689_/X VGND VGND VPWR VPWR _22691_/C sky130_fd_sc_hd__a211o_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21641_ _21250_/X _21640_/X _23914_/Q _21250_/X VGND VGND VPWR VPWR _21641_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21572_ _24097_/Q _21572_/B VGND VGND VPWR VPWR _21572_/X sky130_fd_sc_hd__or2_4
X_24360_ _24361_/CLK _16002_/X HRESETn VGND VGND VPWR VPWR _24360_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20523_ _20522_/X VGND VGND VPWR VPWR _20523_/Y sky130_fd_sc_hd__inv_2
X_23311_ _23135_/CLK _23311_/D VGND VGND VPWR VPWR _23311_/Q sky130_fd_sc_hd__dfxtp_4
X_24291_ _24590_/CLK _24291_/D HRESETn VGND VGND VPWR VPWR _21293_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12564__A _12555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23988__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20454_ _13506_/D _20453_/B _20453_/Y VGND VGND VPWR VPWR _20454_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_119_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23242_ _23242_/CLK _23242_/D VGND VGND VPWR VPWR _19698_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__23917__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20781__A _20800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15875__A _24408_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23173_ _23154_/CLK _19888_/X VGND VGND VPWR VPWR _19887_/A sky130_fd_sc_hd__dfxtp_4
X_20385_ _20385_/A _20385_/B VGND VGND VPWR VPWR _20386_/B sky130_fd_sc_hd__nand2_4
XFILLER_101_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22124_ _21178_/A _22123_/X _21981_/X _15889_/A _16393_/D VGND VGND VPWR VPWR _22124_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_136_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22568__A2 _22011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22055_ _21008_/A VGND VGND VPWR VPWR _22055_/X sky130_fd_sc_hd__buf_2
X_21006_ _21006_/A _19797_/Y VGND VGND VPWR VPWR _21006_/X sky130_fd_sc_hd__or2_4
XFILLER_43_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22501__A _22501_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24776__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21117__A _13324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24705__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22957_ _24496_/Q _22957_/B VGND VGND VPWR VPWR _22957_/X sky130_fd_sc_hd__and2_4
XFILLER_83_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12710_ _12587_/Y _12607_/Y _12554_/X _12710_/D VGND VGND VPWR VPWR _12716_/B sky130_fd_sc_hd__or4_4
XANTENNA__11643__A _11643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22740__A2 _22173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21908_ _17629_/B VGND VGND VPWR VPWR _21924_/A sky130_fd_sc_hd__buf_2
X_13690_ _20201_/B _13687_/X _13688_/Y _13689_/X VGND VGND VPWR VPWR _13691_/B sky130_fd_sc_hd__o22a_4
XFILLER_44_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22888_ _24494_/Q _20757_/A VGND VGND VPWR VPWR _22888_/X sky130_fd_sc_hd__or2_4
XFILLER_70_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12641_ _12578_/Y _12669_/A VGND VGND VPWR VPWR _12641_/X sky130_fd_sc_hd__or2_4
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24627_ _23676_/CLK _15287_/X HRESETn VGND VGND VPWR VPWR _15284_/A sky130_fd_sc_hd__dfstp_4
X_21839_ _21839_/A _11516_/B VGND VGND VPWR VPWR _21839_/X sky130_fd_sc_hd__or2_4
XANTENNA__16965__A2_N _17041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15360_ _22587_/A _15353_/X _11570_/X _15359_/X VGND VGND VPWR VPWR _15360_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_70_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ _24526_/Q VGND VGND VPWR VPWR _12572_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24558_ _24545_/CLK _24558_/D HRESETn VGND VGND VPWR VPWR _24558_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14311_ _20185_/A _14309_/X _20167_/A VGND VGND VPWR VPWR _14311_/X sky130_fd_sc_hd__o21a_4
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11523_ _11496_/Y _11521_/X _11522_/X _11521_/X VGND VGND VPWR VPWR _25220_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23509_ _23514_/CLK _18948_/X VGND VGND VPWR VPWR _17761_/B sky130_fd_sc_hd__dfxtp_4
X_15291_ _14218_/A VGND VGND VPWR VPWR _15291_/X sky130_fd_sc_hd__buf_2
XFILLER_8_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12474__A _12412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24489_ _25090_/CLK _15676_/X HRESETn VGND VGND VPWR VPWR _22736_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17030_ _24030_/Q VGND VGND VPWR VPWR _17030_/Y sky130_fd_sc_hd__inv_2
X_14242_ _14241_/Y _14237_/X _14221_/X _14237_/X VGND VGND VPWR VPWR _14242_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14733__A2 _14732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23658__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14173_ _14172_/X VGND VGND VPWR VPWR _14173_/Y sky130_fd_sc_hd__inv_2
X_13124_ _13230_/A _23132_/Q VGND VGND VPWR VPWR _13125_/C sky130_fd_sc_hd__or2_4
XFILLER_98_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18981_ _18981_/A VGND VGND VPWR VPWR _18981_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15694__B1 _24478_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22114__C _22114_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13055_ _13054_/X VGND VGND VPWR VPWR _13057_/A sky130_fd_sc_hd__inv_2
X_17932_ _17796_/X _18915_/A VGND VGND VPWR VPWR _17933_/C sky130_fd_sc_hd__or2_4
X_12006_ _25140_/Q VGND VGND VPWR VPWR _12006_/Y sky130_fd_sc_hd__inv_2
X_17863_ _17895_/A _23458_/Q VGND VGND VPWR VPWR _17865_/B sky130_fd_sc_hd__or2_4
XFILLER_6_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22411__A _22407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17986__A2 _15430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19602_ _23276_/Q VGND VGND VPWR VPWR _19602_/Y sky130_fd_sc_hd__inv_2
X_16814_ _17067_/A VGND VGND VPWR VPWR _16940_/A sky130_fd_sc_hd__buf_2
X_17794_ _17898_/A _17794_/B _17793_/X VGND VGND VPWR VPWR _17803_/B sky130_fd_sc_hd__or3_4
XANTENNA__22130__B _22524_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16745_ _16745_/A _16731_/X _16739_/X _16745_/D VGND VGND VPWR VPWR _16745_/X sky130_fd_sc_hd__or4_4
X_19533_ _19533_/A VGND VGND VPWR VPWR _19533_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24446__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13957_ _13959_/A _13954_/X _13955_/Y _13956_/X VGND VGND VPWR VPWR _13957_/X sky130_fd_sc_hd__o22a_4
XFILLER_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12908_ _22900_/A _12908_/B VGND VGND VPWR VPWR _12910_/B sky130_fd_sc_hd__or2_4
X_19464_ _19464_/A VGND VGND VPWR VPWR _20993_/B sky130_fd_sc_hd__inv_2
X_16676_ _14592_/B _16023_/X _14589_/B _16024_/Y VGND VGND VPWR VPWR _16680_/C sky130_fd_sc_hd__o22a_4
X_13888_ _13833_/A _13884_/X _13887_/X VGND VGND VPWR VPWR _24912_/D sky130_fd_sc_hd__o21ai_4
XANTENNA__20866__A _20866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15627_ _12546_/Y _15624_/X _15390_/X _15624_/X VGND VGND VPWR VPWR _15627_/X sky130_fd_sc_hd__a2bb2o_4
X_18415_ _18479_/A VGND VGND VPWR VPWR _18469_/A sky130_fd_sc_hd__inv_2
X_12839_ _12838_/Y _24452_/Q _12838_/Y _24452_/Q VGND VGND VPWR VPWR _12844_/B sky130_fd_sc_hd__a2bb2o_4
X_19395_ _18068_/X _11746_/Y _19303_/A _18690_/B VGND VGND VPWR VPWR _19396_/A sky130_fd_sc_hd__or4_4
XFILLER_72_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18346_ _16411_/Y _18472_/A _16411_/Y _23838_/Q VGND VGND VPWR VPWR _18347_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15558_ _15558_/A VGND VGND VPWR VPWR _15558_/X sky130_fd_sc_hd__buf_2
XFILLER_128_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14509_ _24749_/Q _14484_/X _14508_/X VGND VGND VPWR VPWR _14509_/X sky130_fd_sc_hd__a21o_4
X_18277_ _18202_/Y _18277_/B VGND VGND VPWR VPWR _18277_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_171_0_HCLK clkbuf_7_85_0_HCLK/X VGND VGND VPWR VPWR _23282_/CLK sky130_fd_sc_hd__clkbuf_1
X_15489_ _12146_/Y _15487_/X _11563_/X _15487_/X VGND VGND VPWR VPWR _24565_/D sky130_fd_sc_hd__a2bb2o_4
X_17228_ _17228_/A VGND VGND VPWR VPWR _17228_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22247__A1 _23025_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22247__B2 _20866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_28_0_HCLK clkbuf_8_29_0_HCLK/A VGND VGND VPWR VPWR _23925_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12196__C1 _12195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11538__A2 _11535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22798__A2 _22794_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17159_ _17032_/D _17053_/A VGND VGND VPWR VPWR _17160_/B sky130_fd_sc_hd__or2_4
XFILLER_89_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20170_ _23777_/Q _20171_/B VGND VGND VPWR VPWR _20194_/A sky130_fd_sc_hd__and2_4
XFILLER_104_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11728__A _11507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14753__A2_N _14751_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17415__A _17415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23860_ _23762_/CLK _18287_/X HRESETn VGND VGND VPWR VPWR _23860_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24187__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22811_ _21561_/X _22809_/X _21562_/X _22810_/X VGND VGND VPWR VPWR _22811_/X sky130_fd_sc_hd__o22a_4
XFILLER_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23791_ _25183_/CLK MSI_S2 HRESETn VGND VGND VPWR VPWR _23791_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22975__B _23008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24116__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22742_ _22742_/A VGND VGND VPWR VPWR _22743_/C sky130_fd_sc_hd__inv_2
XANTENNA__20776__A _22438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22673_ _22730_/A _22673_/B VGND VGND VPWR VPWR _22687_/C sky130_fd_sc_hd__nor2_4
XFILLER_55_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24412_ _24412_/CLK _15865_/X HRESETn VGND VGND VPWR VPWR _24412_/Q sky130_fd_sc_hd__dfrtp_4
X_21624_ _21612_/A _21624_/B VGND VGND VPWR VPWR _21624_/X sky130_fd_sc_hd__or2_4
XFILLER_90_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24343_ _23872_/CLK _16077_/X HRESETn VGND VGND VPWR VPWR _16075_/A sky130_fd_sc_hd__dfrtp_4
X_21555_ _24918_/Q _22227_/B VGND VGND VPWR VPWR _21555_/X sky130_fd_sc_hd__and2_4
XANTENNA__15699__A1_N _12329_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20506_ _20506_/A VGND VGND VPWR VPWR _20506_/Y sky130_fd_sc_hd__inv_2
X_21486_ _21130_/X _21484_/X _21485_/X VGND VGND VPWR VPWR _21486_/X sky130_fd_sc_hd__and3_4
XFILLER_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23751__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24274_ _24681_/CLK _16263_/X HRESETn VGND VGND VPWR VPWR _24274_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22789__A2 _21562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20437_ _20416_/A VGND VGND VPWR VPWR _20437_/X sky130_fd_sc_hd__buf_2
XANTENNA__21400__A _21400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23225_ _23401_/CLK _19751_/X VGND VGND VPWR VPWR _19749_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_101_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20368_ _20368_/A _20368_/B VGND VGND VPWR VPWR _20369_/B sky130_fd_sc_hd__nand2_4
XANTENNA__18862__B1 _18817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17003__A2_N _24042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23156_ _23156_/CLK _23156_/D VGND VGND VPWR VPWR _23156_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15676__B1 _11558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22107_ _20961_/A _22107_/B VGND VGND VPWR VPWR _22107_/X sky130_fd_sc_hd__or2_4
XANTENNA__11638__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24957__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23087_ _23288_/CLK _20113_/X VGND VGND VPWR VPWR _23087_/Q sky130_fd_sc_hd__dfxtp_4
X_20299_ _14223_/Y _20296_/X _20287_/X _20298_/X VGND VGND VPWR VPWR _20300_/A sky130_fd_sc_hd__a211o_4
XANTENNA__21749__B1 _16393_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22038_ _14045_/Y _11961_/X _15270_/A _20866_/A VGND VGND VPWR VPWR _22038_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22410__A1 _22322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15691__A3 _15505_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22961__A2 _22011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14860_ _24145_/Q VGND VGND VPWR VPWR _14860_/Y sky130_fd_sc_hd__inv_2
X_13811_ _13811_/A _13811_/B _13811_/C _13810_/X VGND VGND VPWR VPWR _13811_/X sky130_fd_sc_hd__and4_4
XFILLER_5_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14791_ _14870_/A VGND VGND VPWR VPWR _14791_/X sky130_fd_sc_hd__buf_2
XFILLER_112_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23989_ _24005_/CLK _17417_/X HRESETn VGND VGND VPWR VPWR _17319_/A sky130_fd_sc_hd__dfrtp_4
X_16530_ _16530_/A VGND VGND VPWR VPWR _16530_/X sky130_fd_sc_hd__buf_2
XFILLER_113_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13742_ _24649_/Q _13742_/B _13742_/C _13742_/D VGND VGND VPWR VPWR _13743_/A sky130_fd_sc_hd__or4_4
XFILLER_44_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23062__A _20740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16461_ _16459_/Y _16460_/X _16373_/X _16460_/X VGND VGND VPWR VPWR _16461_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13673_ _13446_/Y _13671_/X _13638_/X _13671_/X VGND VGND VPWR VPWR _24927_/D sky130_fd_sc_hd__a2bb2o_4
X_18200_ _18256_/A VGND VGND VPWR VPWR _18200_/Y sky130_fd_sc_hd__inv_2
X_15412_ _14020_/A _15314_/X VGND VGND VPWR VPWR _15413_/A sky130_fd_sc_hd__or2_4
XANTENNA__17060__A _17067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12624_ _12629_/A _24505_/Q _12650_/A _12595_/Y VGND VGND VPWR VPWR _12624_/X sky130_fd_sc_hd__a2bb2o_4
X_19180_ _19179_/Y _19175_/X _19089_/X _19175_/X VGND VGND VPWR VPWR _19180_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16392_ _21047_/A VGND VGND VPWR VPWR _16393_/D sky130_fd_sc_hd__buf_2
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23839__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18131_ _18130_/Y _17052_/A _24321_/Q VGND VGND VPWR VPWR _23877_/D sky130_fd_sc_hd__a21oi_4
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15343_ _15342_/Y _15340_/X _11552_/X _15340_/X VGND VGND VPWR VPWR _15343_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12555_ _12554_/X _24518_/Q _12553_/Y _24518_/Q VGND VGND VPWR VPWR _12555_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_244_0_HCLK clkbuf_8_245_0_HCLK/A VGND VGND VPWR VPWR _24264_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11506_ _23763_/Q VGND VGND VPWR VPWR _20842_/B sky130_fd_sc_hd__inv_2
X_18062_ _17459_/Y _18061_/X _17453_/X VGND VGND VPWR VPWR _18062_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__22229__A1 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15274_ _14639_/Y _15272_/X _14232_/X _15272_/X VGND VGND VPWR VPWR _24631_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22229__B2 _22228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12486_ _12465_/B _12464_/X VGND VGND VPWR VPWR _12489_/B sky130_fd_sc_hd__or2_4
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22406__A _16559_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17013_ _16210_/Y _24030_/Q _21124_/A _17160_/A VGND VGND VPWR VPWR _17017_/A sky130_fd_sc_hd__a2bb2o_4
X_14225_ _14047_/A _18633_/A VGND VGND VPWR VPWR _14226_/A sky130_fd_sc_hd__nor2_4
XANTENNA__17105__B1 _17057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21988__B1 _15892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14156_ _12049_/A _12053_/A _14155_/X VGND VGND VPWR VPWR _14156_/X sky130_fd_sc_hd__and3_4
XANTENNA__15667__B1 _11525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13107_ _13102_/X _13104_/X _13106_/X VGND VGND VPWR VPWR _13107_/X sky130_fd_sc_hd__and3_4
XANTENNA__11548__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24698__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14087_ _14086_/Y _14084_/X _13632_/X _14084_/X VGND VGND VPWR VPWR _24859_/D sky130_fd_sc_hd__a2bb2o_4
X_18964_ _18711_/X VGND VGND VPWR VPWR _18964_/X sky130_fd_sc_hd__buf_2
XFILLER_26_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13038_ _11743_/A _13038_/B VGND VGND VPWR VPWR _13038_/X sky130_fd_sc_hd__or2_4
X_17915_ _17947_/A _17911_/X _17915_/C VGND VGND VPWR VPWR _17923_/B sky130_fd_sc_hd__or3_4
X_18895_ _18895_/A VGND VGND VPWR VPWR _18895_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14859__A _14859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19154__A2_N _19146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17846_ _17878_/A _17846_/B VGND VGND VPWR VPWR _17846_/X sky130_fd_sc_hd__or2_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15434__A3 _15432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24280__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14989_ _24711_/Q _14989_/B VGND VGND VPWR VPWR _14989_/X sky130_fd_sc_hd__or2_4
X_17777_ _17815_/A _17777_/B _17777_/C VGND VGND VPWR VPWR _17785_/B sky130_fd_sc_hd__or3_4
XFILLER_47_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19516_ _19510_/Y VGND VGND VPWR VPWR _19516_/X sky130_fd_sc_hd__buf_2
XANTENNA__19030__B1 _18662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16728_ _15943_/Y _17481_/A _15943_/Y _17481_/A VGND VGND VPWR VPWR _16728_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16659_ _16643_/A VGND VGND VPWR VPWR _16659_/X sky130_fd_sc_hd__buf_2
X_19447_ _19447_/A VGND VGND VPWR VPWR _19447_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_54_0_HCLK clkbuf_6_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_54_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19378_ _19372_/Y VGND VGND VPWR VPWR _19378_/X sky130_fd_sc_hd__buf_2
X_18329_ _18300_/A _18327_/X VGND VGND VPWR VPWR _18329_/X sky130_fd_sc_hd__or2_4
X_21340_ _21340_/A _20109_/Y VGND VGND VPWR VPWR _21343_/B sky130_fd_sc_hd__or2_4
XANTENNA__13003__A _12818_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16698__A2 _23960_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21691__A2 _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21271_ _21040_/X _21268_/Y _22245_/A _21270_/X VGND VGND VPWR VPWR _21271_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15370__A2 _15319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16314__A _16339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20222_ _20216_/Y _20221_/X _20209_/A _13711_/X VGND VGND VPWR VPWR _20222_/X sky130_fd_sc_hd__a211o_4
X_23010_ _21546_/X _23007_/Y _22423_/X _23009_/X VGND VGND VPWR VPWR _23010_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20153_ _20152_/Y _20148_/X _15416_/X _20141_/A VGND VGND VPWR VPWR _23069_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24368__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20084_ _23098_/Q VGND VGND VPWR VPWR _20084_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15673__A3 _15596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24961_ _24962_/CLK _24961_/D HRESETn VGND VGND VPWR VPWR _13566_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_134_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23912_ _24928_/CLK _23912_/D HRESETn VGND VGND VPWR VPWR _23912_/Q sky130_fd_sc_hd__dfrtp_4
X_24892_ _24783_/CLK _13965_/X HRESETn VGND VGND VPWR VPWR _24892_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21890__A _21886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23843_ _23824_/CLK _18451_/Y HRESETn VGND VGND VPWR VPWR _23843_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19360__A _11630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23774_ _23774_/CLK _23774_/D HRESETn VGND VGND VPWR VPWR _20192_/A sky130_fd_sc_hd__dfstp_4
X_20986_ _22089_/A _20982_/X _20983_/X _20984_/X _20985_/X VGND VGND VPWR VPWR _20986_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21903__B1 _23660_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22725_ _21529_/X _22723_/X _13362_/A _22724_/X VGND VGND VPWR VPWR _22725_/X sky130_fd_sc_hd__o22a_4
XFILLER_80_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23932__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22656_ _22656_/A VGND VGND VPWR VPWR _22656_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25156__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21607_ _23938_/Q VGND VGND VPWR VPWR _21612_/A sky130_fd_sc_hd__buf_2
XFILLER_107_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14009__A _14009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22587_ _22587_/A _22587_/B VGND VGND VPWR VPWR _22587_/X sky130_fd_sc_hd__and2_4
X_12340_ _25089_/Q _24486_/Q _12412_/C _12339_/Y VGND VGND VPWR VPWR _12340_/X sky130_fd_sc_hd__o22a_4
X_24326_ _23852_/CLK _16122_/X HRESETn VGND VGND VPWR VPWR _16121_/A sky130_fd_sc_hd__dfrtp_4
X_21538_ _21538_/A _21458_/X _21538_/C _21537_/X VGND VGND VPWR VPWR HRDATA[3] sky130_fd_sc_hd__or4_4
XFILLER_127_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12271_ _12176_/A _12280_/B VGND VGND VPWR VPWR _12278_/B sky130_fd_sc_hd__or2_4
Xclkbuf_8_11_0_HCLK clkbuf_7_5_0_HCLK/X VGND VGND VPWR VPWR _23383_/CLK sky130_fd_sc_hd__clkbuf_1
X_24257_ _24654_/CLK _16292_/X HRESETn VGND VGND VPWR VPWR _24257_/Q sky130_fd_sc_hd__dfrtp_4
X_21469_ _21469_/A _21469_/B VGND VGND VPWR VPWR _21471_/B sky130_fd_sc_hd__or2_4
X_14010_ _14000_/B _14008_/Y _13956_/X _14009_/Y _13959_/A VGND VGND VPWR VPWR _14010_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_8_74_0_HCLK clkbuf_8_75_0_HCLK/A VGND VGND VPWR VPWR _24937_/CLK sky130_fd_sc_hd__clkbuf_1
X_23208_ _23303_/CLK _23208_/D VGND VGND VPWR VPWR _19795_/A sky130_fd_sc_hd__dfxtp_4
X_24188_ _24185_/CLK _24188_/D HRESETn VGND VGND VPWR VPWR _24188_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15649__B1 _24500_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24791__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23139_ _23332_/CLK _19978_/X VGND VGND VPWR VPWR _19977_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22135__A1_N _17595_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15961_ _15987_/A VGND VGND VPWR VPWR _15961_/X sky130_fd_sc_hd__buf_2
XFILLER_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23057__A _20735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24720__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14912_ _24674_/Q VGND VGND VPWR VPWR _15138_/B sky130_fd_sc_hd__inv_2
X_17700_ _14573_/A _23422_/Q VGND VGND VPWR VPWR _17702_/B sky130_fd_sc_hd__or2_4
XANTENNA__24038__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15892_ _15892_/A VGND VGND VPWR VPWR _15892_/Y sky130_fd_sc_hd__inv_2
X_18680_ _18677_/Y _18673_/X _18679_/X _18673_/X VGND VGND VPWR VPWR _18680_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11686__B2 _22215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16074__B1 _15770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14843_ _14736_/X _24144_/Q _14736_/X _24144_/Q VGND VGND VPWR VPWR _14843_/X sky130_fd_sc_hd__a2bb2o_4
X_17631_ _23941_/Q VGND VGND VPWR VPWR _17631_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17562_ _17558_/B _17565_/A VGND VGND VPWR VPWR _17563_/B sky130_fd_sc_hd__or2_4
X_14774_ _24704_/Q VGND VGND VPWR VPWR _14809_/A sky130_fd_sc_hd__inv_2
X_11986_ _16475_/A VGND VGND VPWR VPWR _11986_/X sky130_fd_sc_hd__buf_2
XFILLER_63_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16513_ _24175_/Q VGND VGND VPWR VPWR _16513_/Y sky130_fd_sc_hd__inv_2
X_19301_ _19300_/Y _19296_/X _19256_/X _19283_/Y VGND VGND VPWR VPWR _19301_/X sky130_fd_sc_hd__a2bb2o_4
X_13725_ _13745_/B VGND VGND VPWR VPWR _13725_/Y sky130_fd_sc_hd__inv_2
X_17493_ _22395_/A VGND VGND VPWR VPWR _17581_/A sky130_fd_sc_hd__inv_2
XFILLER_72_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17502__B _17502_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11831__A _11830_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16444_ _16443_/Y _16439_/X _16096_/X _16439_/X VGND VGND VPWR VPWR _16444_/X sky130_fd_sc_hd__a2bb2o_4
X_19232_ _18711_/X VGND VGND VPWR VPWR _19232_/X sky130_fd_sc_hd__buf_2
X_13656_ _13655_/Y _13652_/X _11598_/X _13652_/X VGND VGND VPWR VPWR _13656_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14927__A2 _24257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23673__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12607_ _25054_/Q VGND VGND VPWR VPWR _12607_/Y sky130_fd_sc_hd__inv_2
X_19163_ _19162_/Y _19160_/X _19095_/X _19160_/X VGND VGND VPWR VPWR _19163_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16375_ _16375_/A VGND VGND VPWR VPWR _16375_/Y sky130_fd_sc_hd__inv_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13587_ _13586_/X VGND VGND VPWR VPWR _13587_/X sky130_fd_sc_hd__buf_2
XANTENNA__21122__A1 _20885_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18114_ _18110_/Y _18113_/X _18115_/A _18113_/X VGND VGND VPWR VPWR _18114_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15326_ _15401_/A VGND VGND VPWR VPWR _15353_/A sky130_fd_sc_hd__buf_2
X_12538_ _12322_/A _12538_/B VGND VGND VPWR VPWR _12539_/C sky130_fd_sc_hd__or2_4
X_19094_ _19094_/A VGND VGND VPWR VPWR _19094_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22136__A _21245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15888__B1 _15513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18045_ _21147_/A _18044_/X _21147_/A _18044_/X VGND VGND VPWR VPWR _18045_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21040__A _22637_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15257_ _13716_/C _15247_/X _15256_/X _13769_/B _15254_/X VGND VGND VPWR VPWR _24643_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24879__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12469_ _12469_/A _12469_/B VGND VGND VPWR VPWR _12471_/B sky130_fd_sc_hd__or2_4
XANTENNA__16134__A _15655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14208_ _20193_/C VGND VGND VPWR VPWR _20235_/D sky130_fd_sc_hd__inv_2
X_15188_ _14939_/Y _15188_/B VGND VGND VPWR VPWR _15191_/B sky130_fd_sc_hd__or2_4
X_14139_ _24843_/Q _14120_/B _24842_/Q _14115_/X VGND VGND VPWR VPWR _14139_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19445__A _19445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19996_ _19990_/Y VGND VGND VPWR VPWR _19996_/X sky130_fd_sc_hd__buf_2
XANTENNA__13115__A1 _11711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24461__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18947_ _17761_/B VGND VGND VPWR VPWR _18947_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21189__A1 _22806_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22386__B1 _24515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22925__A2 _22859_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18878_ _18872_/Y _18877_/X _18764_/X _18877_/X VGND VGND VPWR VPWR _18878_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16065__B1 _15761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17829_ _17935_/A _23579_/Q VGND VGND VPWR VPWR _17829_/X sky130_fd_sc_hd__or2_4
X_20840_ _12793_/Y _20837_/X _20839_/X VGND VGND VPWR VPWR _20840_/X sky130_fd_sc_hd__a21o_4
XANTENNA__22689__A1 _14900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20771_ _17032_/D _22201_/A _20748_/X _20770_/X VGND VGND VPWR VPWR _20772_/A sky130_fd_sc_hd__a211o_4
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21361__B2 _22548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22510_ _11949_/A _22510_/B _22510_/C _21033_/X VGND VGND VPWR VPWR _22510_/X sky130_fd_sc_hd__or4_4
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23490_ _23489_/CLK _19001_/X VGND VGND VPWR VPWR _23490_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15040__A1 _15033_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22441_ _21572_/B _22439_/X _22441_/C VGND VGND VPWR VPWR _22441_/X sky130_fd_sc_hd__and3_4
XFILLER_91_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13364__A1_N _11913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25160_ _23885_/CLK _25160_/D HRESETn VGND VGND VPWR VPWR _25160_/Q sky130_fd_sc_hd__dfrtp_4
X_22372_ _22371_/X VGND VGND VPWR VPWR _22372_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22861__A1 _14859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24111_ _24698_/CLK _16645_/X HRESETn VGND VGND VPWR VPWR _14722_/A sky130_fd_sc_hd__dfrtp_4
X_21323_ _21323_/A _21323_/B _21323_/C _21323_/D VGND VGND VPWR VPWR _21323_/X sky130_fd_sc_hd__or4_4
XANTENNA__13668__A _13668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25091_ _25091_/CLK _25091_/D HRESETn VGND VGND VPWR VPWR _12469_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_117_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21254_ _21253_/X VGND VGND VPWR VPWR _21254_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24549__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24042_ _24042_/CLK _24042_/D HRESETn VGND VGND VPWR VPWR _24042_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20205_ _20204_/X VGND VGND VPWR VPWR _20205_/Y sky130_fd_sc_hd__inv_2
X_21185_ _21180_/X _21184_/Y _11677_/Y _21180_/X VGND VGND VPWR VPWR _21185_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19355__A _19349_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20136_ _20141_/A VGND VGND VPWR VPWR _20136_/X sky130_fd_sc_hd__buf_2
XANTENNA__15646__A3 _15635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24131__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20067_ _20060_/A VGND VGND VPWR VPWR _20067_/X sky130_fd_sc_hd__buf_2
XANTENNA__19242__B1 _11839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24944_ _24944_/CLK _24944_/D HRESETn VGND VGND VPWR VPWR _24944_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21109__B _21109_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11668__B2 _22450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22392__A3 _22251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24875_ _23657_/CLK _24875_/D HRESETn VGND VGND VPWR VPWR _24875_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15803__B1 _15709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11840_ _11830_/Y VGND VGND VPWR VPWR _11840_/X sky130_fd_sc_hd__buf_2
X_23826_ _23826_/CLK _23826_/D HRESETn VGND VGND VPWR VPWR _18517_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_96_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11771_ _17448_/B VGND VGND VPWR VPWR _11771_/Y sky130_fd_sc_hd__inv_2
X_23757_ _24185_/CLK _23757_/D HRESETn VGND VGND VPWR VPWR _23757_/Q sky130_fd_sc_hd__dfrtp_4
X_20969_ _20962_/X _20967_/X _20968_/X VGND VGND VPWR VPWR _20969_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12747__A _12749_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16219__A _14218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13510_ _20520_/A _13510_/B _13509_/X VGND VGND VPWR VPWR _13510_/X sky130_fd_sc_hd__or3_4
X_22708_ _22707_/X VGND VGND VPWR VPWR _22708_/Y sky130_fd_sc_hd__inv_2
X_14490_ _14489_/X VGND VGND VPWR VPWR _14490_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16244__A1_N _14920_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23688_ _24879_/CLK _23688_/D HRESETn VGND VGND VPWR VPWR _23688_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13441_ _24925_/Q VGND VGND VPWR VPWR _13441_/Y sky130_fd_sc_hd__inv_2
X_22639_ _22639_/A _22638_/X VGND VGND VPWR VPWR _22639_/X sky130_fd_sc_hd__or2_4
X_16160_ _16160_/A VGND VGND VPWR VPWR _16160_/Y sky130_fd_sc_hd__inv_2
X_13372_ _13363_/A VGND VGND VPWR VPWR _13372_/X sky130_fd_sc_hd__buf_2
X_15111_ _24651_/Q VGND VGND VPWR VPWR _15112_/C sky130_fd_sc_hd__inv_2
XFILLER_6_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12323_ _12405_/D _20808_/A _12405_/D _20808_/A VGND VGND VPWR VPWR _12323_/X sky130_fd_sc_hd__a2bb2o_4
X_24309_ _24604_/CLK _16168_/X HRESETn VGND VGND VPWR VPWR _24309_/Q sky130_fd_sc_hd__dfrtp_4
X_16091_ _16089_/Y _16084_/X _11585_/X _16090_/X VGND VGND VPWR VPWR _24338_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24972__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15042_ _15042_/A _15019_/X VGND VGND VPWR VPWR _15043_/A sky130_fd_sc_hd__or2_4
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12254_ _12254_/A VGND VGND VPWR VPWR _12254_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24901__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19850_ _21669_/B _19847_/X _19825_/X _19847_/X VGND VGND VPWR VPWR _23187_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24219__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12185_ _12185_/A _12185_/B _12184_/X VGND VGND VPWR VPWR _12192_/A sky130_fd_sc_hd__or3_4
XANTENNA__19481__B1 _19387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16295__B1 _16219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18801_ HWDATA[1] VGND VGND VPWR VPWR _18801_/X sky130_fd_sc_hd__buf_2
X_19781_ _19780_/Y VGND VGND VPWR VPWR _19781_/X sky130_fd_sc_hd__buf_2
XFILLER_95_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16993_ _24306_/Q _16992_/Y _16205_/Y _24032_/Q VGND VGND VPWR VPWR _16999_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_135_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18732_ _17678_/B VGND VGND VPWR VPWR _18732_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19233__B1 _19232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15944_ _15943_/Y _15941_/X _11555_/X _15941_/X VGND VGND VPWR VPWR _24383_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16047__B1 _15828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15875_ _24408_/Q VGND VGND VPWR VPWR _15875_/Y sky130_fd_sc_hd__inv_2
X_18663_ _21001_/B _18657_/X _18662_/X _18644_/Y VGND VGND VPWR VPWR _18663_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14826_ _24712_/Q _24155_/Q _14977_/C _14825_/Y VGND VGND VPWR VPWR _14829_/C sky130_fd_sc_hd__o22a_4
X_17614_ _17614_/A _17614_/B VGND VGND VPWR VPWR _17615_/B sky130_fd_sc_hd__or2_4
XFILLER_52_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18594_ _16325_/A _18470_/A _16325_/A _18470_/A VGND VGND VPWR VPWR _18597_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23854__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25078__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21035__A _21034_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14757_ _14757_/A VGND VGND VPWR VPWR _14757_/Y sky130_fd_sc_hd__inv_2
X_17545_ _17528_/X _17545_/B _17544_/X VGND VGND VPWR VPWR _17545_/X sky130_fd_sc_hd__or3_4
XFILLER_75_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11969_ _11968_/Y _11966_/X _11616_/X _11966_/X VGND VGND VPWR VPWR _25154_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12084__B2 _24561_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16129__A _14197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25007__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13708_ _24914_/Q _13686_/X _23126_/Q _13681_/X VGND VGND VPWR VPWR _13708_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15033__A _15033_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17476_ _16746_/X VGND VGND VPWR VPWR _17619_/A sky130_fd_sc_hd__buf_2
X_14688_ _14062_/Y _14621_/X _14647_/X _14687_/Y VGND VGND VPWR VPWR _14689_/A sky130_fd_sc_hd__o22a_4
XFILLER_32_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19215_ _21876_/A VGND VGND VPWR VPWR _19215_/Y sky130_fd_sc_hd__inv_2
X_13639_ _13630_/X VGND VGND VPWR VPWR _13639_/X sky130_fd_sc_hd__buf_2
X_16427_ _16425_/Y _16421_/X _16261_/X _16426_/X VGND VGND VPWR VPWR _24209_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22027__A1_N _13934_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16358_ _16358_/A VGND VGND VPWR VPWR _16358_/Y sky130_fd_sc_hd__inv_2
X_19146_ _19153_/A VGND VGND VPWR VPWR _19146_/X sky130_fd_sc_hd__buf_2
XANTENNA__11595__B1 _11594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15309_ _21300_/A VGND VGND VPWR VPWR _21581_/A sky130_fd_sc_hd__buf_2
X_16289_ _15915_/X _16276_/X _15706_/X _24258_/Q _16237_/A VGND VGND VPWR VPWR _16289_/X
+ sky130_fd_sc_hd__a32o_4
X_19077_ _17677_/B VGND VGND VPWR VPWR _19077_/Y sky130_fd_sc_hd__inv_2
X_18028_ _19531_/A VGND VGND VPWR VPWR _18030_/A sky130_fd_sc_hd__inv_2
XANTENNA__24642__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19979_ _19979_/A VGND VGND VPWR VPWR _21521_/B sky130_fd_sc_hd__inv_2
XFILLER_45_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19224__B1 _19201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22990_ _23023_/A _22990_/B _22990_/C VGND VGND VPWR VPWR _22990_/X sky130_fd_sc_hd__and3_4
XANTENNA__19775__B2 _19772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21941_ _21500_/A _21939_/X _21940_/X VGND VGND VPWR VPWR _21941_/X sky130_fd_sc_hd__and3_4
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20768__B _22445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24660_ _24662_/CLK _15207_/X HRESETn VGND VGND VPWR VPWR _24660_/Q sky130_fd_sc_hd__dfrtp_4
X_21872_ _23084_/Q _15639_/X VGND VGND VPWR VPWR _21872_/X sky130_fd_sc_hd__and2_4
XPHY_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ _23482_/CLK _18653_/X VGND VGND VPWR VPWR _23611_/Q sky130_fd_sc_hd__dfxtp_4
X_20823_ _20802_/X VGND VGND VPWR VPWR _20823_/X sky130_fd_sc_hd__buf_2
XANTENNA__15800__A3 _15706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24591_ _23702_/CLK _24591_/D HRESETn VGND VGND VPWR VPWR _15385_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_78_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22983__B _22857_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23542_ _23133_/CLK _18855_/X VGND VGND VPWR VPWR _13039_/B sky130_fd_sc_hd__dfxtp_4
X_20754_ _15908_/Y _23025_/B VGND VGND VPWR VPWR _20754_/X sky130_fd_sc_hd__or2_4
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23473_ _24998_/CLK _19050_/X VGND VGND VPWR VPWR _23473_/Q sky130_fd_sc_hd__dfxtp_4
X_20685_ _23926_/Q _13474_/A _15810_/B _15807_/A _15720_/X VGND VGND VPWR VPWR _20685_/X
+ sky130_fd_sc_hd__o32a_4
Xclkbuf_5_24_0_HCLK clkbuf_4_12_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_49_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25212_ _25214_/CLK _25212_/D HRESETn VGND VGND VPWR VPWR _25212_/Q sky130_fd_sc_hd__dfrtp_4
X_22424_ _12362_/A _11964_/A VGND VGND VPWR VPWR _22424_/X sky130_fd_sc_hd__or2_4
XFILLER_13_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11586__B1 _11585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13398__A _13398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25143_ _23789_/CLK _25143_/D HRESETn VGND VGND VPWR VPWR _11999_/A sky130_fd_sc_hd__dfrtp_4
X_22355_ _22355_/A _20911_/X VGND VGND VPWR VPWR _22355_/X sky130_fd_sc_hd__and2_4
X_21306_ _21305_/X VGND VGND VPWR VPWR _21323_/B sky130_fd_sc_hd__inv_2
XANTENNA__24383__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25074_ _23716_/CLK _12528_/Y HRESETn VGND VGND VPWR VPWR _21566_/A sky130_fd_sc_hd__dfrtp_4
X_22286_ _23737_/Q _22173_/X _23705_/Q _22285_/X VGND VGND VPWR VPWR _22286_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_85_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24312__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24025_ _23664_/CLK _24025_/D HRESETn VGND VGND VPWR VPWR _24025_/Q sky130_fd_sc_hd__dfstp_4
X_21237_ _21237_/A VGND VGND VPWR VPWR _21394_/A sky130_fd_sc_hd__buf_2
XFILLER_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16277__B1 _22312_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21168_ _17651_/A VGND VGND VPWR VPWR _21169_/A sky130_fd_sc_hd__buf_2
XFILLER_133_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_148_0_HCLK clkbuf_7_74_0_HCLK/X VGND VGND VPWR VPWR _25214_/CLK sky130_fd_sc_hd__clkbuf_1
X_20119_ _22218_/C VGND VGND VPWR VPWR _20119_/X sky130_fd_sc_hd__buf_2
X_13990_ _13956_/X _13989_/X _24812_/Q _13959_/A VGND VGND VPWR VPWR _13990_/Y sky130_fd_sc_hd__a22oi_4
X_21099_ _16300_/A _21098_/X VGND VGND VPWR VPWR _21099_/X sky130_fd_sc_hd__or2_4
XANTENNA__14022__A _14197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12941_ _12854_/Y _12935_/X _12922_/X _12937_/Y VGND VGND VPWR VPWR _12942_/A sky130_fd_sc_hd__a211o_4
X_24927_ _24757_/CLK _24927_/D HRESETn VGND VGND VPWR VPWR _13446_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15660_ _15664_/A VGND VGND VPWR VPWR _15661_/A sky130_fd_sc_hd__buf_2
XFILLER_73_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12872_ _12774_/Y _21840_/A VGND VGND VPWR VPWR _12878_/B sky130_fd_sc_hd__or2_4
XFILLER_18_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24858_ _23657_/CLK _24858_/D HRESETn VGND VGND VPWR VPWR _24858_/Q sky130_fd_sc_hd__dfrtp_4
X_14611_ _24721_/Q _14610_/X _14626_/A VGND VGND VPWR VPWR _14612_/B sky130_fd_sc_hd__or3_4
XANTENNA__25171__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11823_ _11823_/A _11814_/Y VGND VGND VPWR VPWR _11823_/Y sky130_fd_sc_hd__nor2_4
XFILLER_57_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23809_ _23624_/CLK _18627_/X HRESETn VGND VGND VPWR VPWR _23809_/Q sky130_fd_sc_hd__dfstp_4
X_15591_ _12579_/Y _15590_/X _11525_/X _15590_/X VGND VGND VPWR VPWR _24531_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12477__A _12474_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24789_ _24823_/CLK _14294_/X HRESETn VGND VGND VPWR VPWR _24789_/Q sky130_fd_sc_hd__dfrtp_4
X_17330_ _17330_/A _17329_/X VGND VGND VPWR VPWR _17331_/A sky130_fd_sc_hd__or2_4
XANTENNA__25100__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14542_/A _14482_/X VGND VGND VPWR VPWR _14543_/A sky130_fd_sc_hd__or2_4
XPHY_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11757_/A VGND VGND VPWR VPWR _11755_/A sky130_fd_sc_hd__buf_2
XPHY_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16201__B1 _15890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _25219_/Q _24007_/Q _11524_/Y _17260_/Y VGND VGND VPWR VPWR _17261_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15788__A _15788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _14471_/X _14445_/A _21396_/A _14445_/Y VGND VGND VPWR VPWR _14473_/X sky130_fd_sc_hd__o22a_4
XPHY_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _11685_/A VGND VGND VPWR VPWR _13585_/A sky130_fd_sc_hd__inv_2
XFILLER_35_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16752__B2 _16846_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16212_ _16210_/Y _16208_/X _16211_/X _16208_/X VGND VGND VPWR VPWR _16212_/X sky130_fd_sc_hd__a2bb2o_4
X_19000_ _23490_/Q VGND VGND VPWR VPWR _19000_/Y sky130_fd_sc_hd__inv_2
XPHY_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13424_ _13655_/A _14385_/A _24934_/Q _14383_/A VGND VGND VPWR VPWR _13427_/C sky130_fd_sc_hd__a2bb2o_4
X_17192_ _17171_/X _17185_/X _24022_/Q _20723_/A _17188_/X VGND VGND VPWR VPWR _24023_/D
+ sky130_fd_sc_hd__a32o_4
X_16143_ _24318_/Q VGND VGND VPWR VPWR _16143_/Y sky130_fd_sc_hd__inv_2
X_13355_ _24987_/Q VGND VGND VPWR VPWR _13355_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12306_ _12305_/Y _24498_/Q _12305_/Y _24498_/Q VGND VGND VPWR VPWR _12312_/B sky130_fd_sc_hd__a2bb2o_4
X_16074_ _16073_/Y _16071_/X _15770_/X _16071_/X VGND VGND VPWR VPWR _16074_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13286_ _13222_/A _13282_/X _13285_/X VGND VGND VPWR VPWR _13287_/C sky130_fd_sc_hd__or3_4
XFILLER_53_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15025_ _14874_/Y _15025_/B VGND VGND VPWR VPWR _15026_/C sky130_fd_sc_hd__or2_4
X_19902_ _19901_/Y _19897_/X _19859_/X _19897_/A VGND VGND VPWR VPWR _19902_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24053__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12237_ _12237_/A _12228_/X VGND VGND VPWR VPWR _12237_/X sky130_fd_sc_hd__or2_4
XANTENNA__17508__A _23012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_44_0_HCLK clkbuf_7_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_44_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12541__A2 _12434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21261__B1 _21793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19833_ _19830_/Y _19831_/X _19832_/X _19831_/X VGND VGND VPWR VPWR _19833_/X sky130_fd_sc_hd__a2bb2o_4
X_12168_ _12167_/Y VGND VGND VPWR VPWR _12186_/B sky130_fd_sc_hd__buf_2
X_19764_ _19764_/A VGND VGND VPWR VPWR _21812_/B sky130_fd_sc_hd__inv_2
X_12099_ _12097_/A _12098_/A _12097_/Y _12098_/Y VGND VGND VPWR VPWR _12099_/X sky130_fd_sc_hd__o22a_4
X_16976_ _16198_/A _22164_/A _16198_/Y _17145_/A VGND VGND VPWR VPWR _16981_/B sky130_fd_sc_hd__o22a_4
XFILLER_110_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20869__A _14009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18715_ _18714_/Y _14594_/X _17199_/X _14594_/X VGND VGND VPWR VPWR _23590_/D sky130_fd_sc_hd__a2bb2o_4
X_15927_ _24389_/Q VGND VGND VPWR VPWR _15927_/Y sky130_fd_sc_hd__inv_2
X_19695_ _19693_/Y _19689_/X _19603_/X _19694_/X VGND VGND VPWR VPWR _19695_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22761__B1 _24525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18646_ _22056_/B _18645_/X _15541_/X _18645_/X VGND VGND VPWR VPWR _23614_/D sky130_fd_sc_hd__a2bb2o_4
X_15858_ _15857_/Y _15854_/X _15770_/X _15854_/X VGND VGND VPWR VPWR _24415_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16440__B1 _15369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14809_ _14809_/A VGND VGND VPWR VPWR _15003_/A sky130_fd_sc_hd__buf_2
XFILLER_18_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12057__A1 _12011_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18577_ _16363_/A _23822_/Q _16363_/Y _18532_/A VGND VGND VPWR VPWR _18577_/X sky130_fd_sc_hd__o22a_4
X_15789_ _12787_/Y _15787_/X _15788_/X _15787_/X VGND VGND VPWR VPWR _15789_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17528_ _16747_/Y VGND VGND VPWR VPWR _17528_/X sky130_fd_sc_hd__buf_2
XANTENNA__24894__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17459_ _21491_/A VGND VGND VPWR VPWR _17459_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24823__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20470_ _20468_/Y _20462_/Y _20469_/X VGND VGND VPWR VPWR _20470_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16306__B _16306_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19129_ _17772_/B VGND VGND VPWR VPWR _19129_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22140_ _11904_/Y _14013_/B _21581_/A VGND VGND VPWR VPWR _22140_/X sky130_fd_sc_hd__o21a_4
XFILLER_134_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22071_ _22055_/X _22071_/B VGND VGND VPWR VPWR _22071_/X sky130_fd_sc_hd__or2_4
XFILLER_133_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17418__A _17415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22043__B _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21022_ _13526_/B _21069_/A VGND VGND VPWR VPWR _21022_/X sky130_fd_sc_hd__and2_4
XANTENNA__16274__A3 _16093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23776__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_1_0_HCLK clkbuf_6_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_75_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20779__A _22933_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19748__B2 _19743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20874__A2_N _21590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23705__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22973_ _23026_/B _22972_/X _22459_/X _24532_/Q _22460_/X VGND VGND VPWR VPWR _22974_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14777__A _14777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17153__A _17129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24712_ _24712_/CLK _14986_/Y HRESETn VGND VGND VPWR VPWR _24712_/Q sky130_fd_sc_hd__dfrtp_4
X_21924_ _21924_/A _19691_/Y VGND VGND VPWR VPWR _21924_/X sky130_fd_sc_hd__or2_4
XFILLER_56_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16431__B1 _16266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24815__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24643_ _24643_/CLK _24643_/D HRESETn VGND VGND VPWR VPWR _13716_/B sky130_fd_sc_hd__dfrtp_4
X_21855_ _21256_/X _21855_/B _21855_/C _21855_/D VGND VGND VPWR VPWR _21855_/X sky130_fd_sc_hd__or4_4
XFILLER_70_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ _20806_/A VGND VGND VPWR VPWR _20832_/A sky130_fd_sc_hd__buf_2
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24574_ _24545_/CLK _15473_/X HRESETn VGND VGND VPWR VPWR _24574_/Q sky130_fd_sc_hd__dfrtp_4
X_21786_ _21786_/A _21786_/B VGND VGND VPWR VPWR _21786_/X sky130_fd_sc_hd__or2_4
XANTENNA__18184__B1 _16073_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23525_ _23531_/CLK _23525_/D VGND VGND VPWR VPWR _17757_/B sky130_fd_sc_hd__dfxtp_4
X_20737_ _20737_/A _20737_/B VGND VGND VPWR VPWR _20737_/X sky130_fd_sc_hd__and2_4
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22218__B _22024_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13548__A1 _20883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15401__A _15401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22807__A1 _16061_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24564__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23456_ _23568_/CLK _23456_/D VGND VGND VPWR VPWR _19094_/A sky130_fd_sc_hd__dfxtp_4
X_20668_ _20647_/X _20667_/Y _24184_/Q _20651_/X VGND VGND VPWR VPWR _20668_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22407_ _22407_/A VGND VGND VPWR VPWR _22407_/X sky130_fd_sc_hd__buf_2
XANTENNA__11627__A1_N _11623_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19808__A _11635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23387_ _23388_/CLK _23387_/D VGND VGND VPWR VPWR _23387_/Q sky130_fd_sc_hd__dfxtp_4
X_20599_ _20599_/A VGND VGND VPWR VPWR _20599_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18712__A _18711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20294__A1 _14230_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13140_ _13244_/A _13140_/B VGND VGND VPWR VPWR _13142_/B sky130_fd_sc_hd__or2_4
X_25126_ _25130_/CLK _25126_/D HRESETn VGND VGND VPWR VPWR _25126_/Q sky130_fd_sc_hd__dfrtp_4
X_22338_ _22338_/A VGND VGND VPWR VPWR _22338_/X sky130_fd_sc_hd__buf_2
XFILLER_100_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13071_ _13230_/A _23133_/Q VGND VGND VPWR VPWR _13072_/C sky130_fd_sc_hd__or2_4
X_25057_ _24523_/CLK _12707_/Y HRESETn VGND VGND VPWR VPWR _25057_/Q sky130_fd_sc_hd__dfrtp_4
X_22269_ _22225_/X _22266_/X _22231_/X _22268_/X VGND VGND VPWR VPWR _22270_/B sky130_fd_sc_hd__o22a_4
XANTENNA__16232__A _16235_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12022_ _12022_/A VGND VGND VPWR VPWR _12022_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21243__B1 _21242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24008_ _24008_/CLK _17338_/Y HRESETn VGND VGND VPWR VPWR _24008_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17998__B1 _23914_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22888__B _20757_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16830_ _24071_/Q VGND VGND VPWR VPWR _16839_/B sky130_fd_sc_hd__inv_2
XANTENNA__16670__B1 _24096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19739__B2 _19738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13973_ _13959_/A VGND VGND VPWR VPWR _13973_/X sky130_fd_sc_hd__buf_2
X_16761_ _24086_/Q VGND VGND VPWR VPWR _16866_/A sky130_fd_sc_hd__inv_2
XFILLER_58_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18500_ _18358_/Y _18504_/B VGND VGND VPWR VPWR _18501_/C sky130_fd_sc_hd__nand2_4
XFILLER_46_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12924_ _12923_/X VGND VGND VPWR VPWR _12924_/Y sky130_fd_sc_hd__inv_2
X_15712_ _15712_/A VGND VGND VPWR VPWR _15712_/X sky130_fd_sc_hd__buf_2
XFILLER_59_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16692_ _16692_/A VGND VGND VPWR VPWR _16692_/Y sky130_fd_sc_hd__inv_2
X_19480_ _19467_/Y VGND VGND VPWR VPWR _19480_/X sky130_fd_sc_hd__buf_2
XFILLER_92_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16422__B1 _16334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18431_ _23827_/Q VGND VGND VPWR VPWR _18486_/B sky130_fd_sc_hd__inv_2
XFILLER_98_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12855_ _12845_/A _12853_/Y _12854_/Y _24449_/Q VGND VGND VPWR VPWR _12855_/X sky130_fd_sc_hd__a2bb2o_4
X_15643_ _15642_/X VGND VGND VPWR VPWR _21795_/B sky130_fd_sc_hd__buf_2
X_11806_ _11809_/B _11804_/A _11815_/C _11805_/X VGND VGND VPWR VPWR _11807_/A sky130_fd_sc_hd__o22a_4
X_15574_ _16624_/A VGND VGND VPWR VPWR _15574_/X sky130_fd_sc_hd__buf_2
X_18362_ _24198_/Q _23821_/Q _16454_/Y _18536_/A VGND VGND VPWR VPWR _18362_/X sky130_fd_sc_hd__o22a_4
X_12786_ _12943_/C _24445_/Q _12943_/C _24445_/Q VGND VGND VPWR VPWR _12795_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18175__B1 _24345_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14471_/X _14524_/X _14471_/X _14524_/X VGND VGND VPWR VPWR _24746_/D sky130_fd_sc_hd__a2bb2o_4
X_17313_ _17266_/Y _17270_/Y _17312_/X VGND VGND VPWR VPWR _17313_/X sky130_fd_sc_hd__or3_4
XPHY_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11737_ _11733_/X VGND VGND VPWR VPWR _11737_/Y sky130_fd_sc_hd__inv_2
XPHY_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18293_ _18295_/B VGND VGND VPWR VPWR _18294_/B sky130_fd_sc_hd__inv_2
XANTENNA__15528__A2 _15319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16725__B2 _22434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14456_ _21237_/A VGND VGND VPWR VPWR _14524_/A sky130_fd_sc_hd__buf_2
X_17244_ _17244_/A VGND VGND VPWR VPWR _17415_/A sky130_fd_sc_hd__inv_2
XANTENNA__21032__B _21408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11668_ _11667_/Y _22450_/A _11667_/Y _22450_/A VGND VGND VPWR VPWR _11668_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _13407_/A _13407_/B VGND VGND VPWR VPWR _13456_/A sky130_fd_sc_hd__and2_4
XANTENNA__20809__B1 _20807_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17175_ _23671_/Q _17174_/X VGND VGND VPWR VPWR _20368_/B sky130_fd_sc_hd__or2_4
XANTENNA__15030__B _15034_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24234__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14387_ _14387_/A _14386_/Y _14387_/C _24767_/Q VGND VGND VPWR VPWR _14387_/X sky130_fd_sc_hd__and4_4
X_11599_ _11599_/A VGND VGND VPWR VPWR _11599_/X sky130_fd_sc_hd__buf_2
XFILLER_128_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16126_ _16125_/Y _16046_/A _15291_/X _16046_/A VGND VGND VPWR VPWR _24324_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_6_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16489__B1 _16246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13338_ _14047_/A _13328_/X VGND VGND VPWR VPWR _13338_/Y sky130_fd_sc_hd__nor2_4
XFILLER_109_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16057_ _16056_/Y _16052_/X _15756_/X _16052_/X VGND VGND VPWR VPWR _24351_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13269_ _13301_/A _13269_/B VGND VGND VPWR VPWR _13270_/C sky130_fd_sc_hd__or2_4
X_15008_ _14703_/X _15006_/A VGND VGND VPWR VPWR _15008_/X sky130_fd_sc_hd__or2_4
XANTENNA__20037__B2 _20036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17989__B1 _15788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19816_ _22072_/B _19814_/X _19815_/X _19814_/X VGND VGND VPWR VPWR _19816_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25093__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_131_0_HCLK clkbuf_7_65_0_HCLK/X VGND VGND VPWR VPWR _23469_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_96_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16661__B1 _15788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19747_ _19747_/A VGND VGND VPWR VPWR _21482_/B sky130_fd_sc_hd__inv_2
X_16959_ _16190_/Y _24038_/Q _16190_/Y _24038_/Q VGND VGND VPWR VPWR _16959_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21537__A1 _21530_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_194_0_HCLK clkbuf_7_97_0_HCLK/X VGND VGND VPWR VPWR _24319_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25022__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19678_ _19677_/Y _19673_/X _19610_/X _19673_/X VGND VGND VPWR VPWR _23250_/D sky130_fd_sc_hd__a2bb2o_4
X_18629_ _18607_/X _18621_/X _20705_/B _23807_/Q _18624_/X VGND VGND VPWR VPWR _18629_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_53_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22901__A2_N _22178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13006__A _12925_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21640_ _20892_/X _21639_/X _18005_/Y _22616_/A VGND VGND VPWR VPWR _21640_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21223__A _21383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21571_ _21298_/B VGND VGND VPWR VPWR _21572_/B sky130_fd_sc_hd__buf_2
XFILLER_20_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23310_ _23308_/CLK _19512_/X VGND VGND VPWR VPWR _23310_/Q sky130_fd_sc_hd__dfxtp_4
X_20522_ _22753_/A _20416_/A _20446_/X _20521_/X VGND VGND VPWR VPWR _20522_/X sky130_fd_sc_hd__o22a_4
X_24290_ _24289_/CLK _16217_/X HRESETn VGND VGND VPWR VPWR _21124_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23241_ _23385_/CLK _23241_/D VGND VGND VPWR VPWR _23241_/Q sky130_fd_sc_hd__dfxtp_4
X_20453_ _13506_/D _20453_/B VGND VGND VPWR VPWR _20453_/Y sky130_fd_sc_hd__nor2_4
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23172_ _23332_/CLK _23172_/D VGND VGND VPWR VPWR _23172_/Q sky130_fd_sc_hd__dfxtp_4
X_20384_ _20383_/X VGND VGND VPWR VPWR _20384_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22123_ _16200_/A _21979_/X VGND VGND VPWR VPWR _22123_/X sky130_fd_sc_hd__or2_4
XFILLER_97_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21557__A2_N _21178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23957__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20028__B2 _20027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22054_ _21665_/A _22052_/X _22053_/X VGND VGND VPWR VPWR _22059_/B sky130_fd_sc_hd__and3_4
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22973__B1 _24532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21005_ _20998_/A _19986_/Y VGND VGND VPWR VPWR _21005_/X sky130_fd_sc_hd__or2_4
XANTENNA__19363__A _19349_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17444__A2 _17366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_90_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_90_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22725__B1 _13362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22956_ _12432_/A _22956_/B VGND VGND VPWR VPWR _22956_/X sky130_fd_sc_hd__or2_4
XFILLER_83_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21907_ _22223_/A _21885_/X _21890_/Y _21895_/X _21906_/X VGND VGND VPWR VPWR _21907_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_56_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22887_ _22931_/A _22880_/X _22882_/X _22585_/A _22886_/Y VGND VGND VPWR VPWR _22887_/X
+ sky130_fd_sc_hd__a32o_4
X_12640_ _25065_/Q VGND VGND VPWR VPWR _12669_/A sky130_fd_sc_hd__inv_2
XFILLER_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24626_ _24870_/CLK _24626_/D HRESETn VGND VGND VPWR VPWR _15288_/A sky130_fd_sc_hd__dfstp_4
X_21838_ _21837_/X VGND VGND VPWR VPWR _21838_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24745__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21133__A _21153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ _25061_/Q VGND VGND VPWR VPWR _12571_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24557_ _24545_/CLK _24557_/D HRESETn VGND VGND VPWR VPWR _24557_/Q sky130_fd_sc_hd__dfrtp_4
X_21769_ _21760_/X _21769_/B VGND VGND VPWR VPWR _21769_/X sky130_fd_sc_hd__or2_4
XFILLER_93_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14310_ _13863_/A _20175_/A VGND VGND VPWR VPWR _20167_/A sky130_fd_sc_hd__or2_4
XFILLER_19_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11522_ HWDATA[30] VGND VGND VPWR VPWR _11522_/X sky130_fd_sc_hd__buf_2
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23508_ _23514_/CLK _23508_/D VGND VGND VPWR VPWR _18949_/A sky130_fd_sc_hd__dfxtp_4
X_15290_ _15290_/A VGND VGND VPWR VPWR _15290_/Y sky130_fd_sc_hd__inv_2
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24488_ _24488_/CLK _15678_/X HRESETn VGND VGND VPWR VPWR _24488_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20972__A _20972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14241_ _24811_/Q VGND VGND VPWR VPWR _14241_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15391__B1 _15390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23439_ _23440_/CLK _23439_/D VGND VGND VPWR VPWR _23439_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_109_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14172_ _14159_/Y _14155_/X _14145_/X _14171_/X VGND VGND VPWR VPWR _14172_/X sky130_fd_sc_hd__a211o_4
X_13123_ _13300_/A _13123_/B VGND VGND VPWR VPWR _13125_/B sky130_fd_sc_hd__or2_4
X_25109_ _25115_/CLK _25109_/D HRESETn VGND VGND VPWR VPWR _25109_/Q sky130_fd_sc_hd__dfrtp_4
X_18980_ _18979_/Y _18975_/X _18932_/X _18975_/X VGND VGND VPWR VPWR _23498_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23698__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13054_ _11868_/Y _13053_/X _11871_/C VGND VGND VPWR VPWR _13054_/X sky130_fd_sc_hd__o21a_4
X_17931_ _17899_/A _18893_/A VGND VGND VPWR VPWR _17931_/X sky130_fd_sc_hd__or2_4
XANTENNA__22114__D _22113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12005_ _12004_/Y _12002_/X _11631_/X _12002_/X VGND VGND VPWR VPWR _25141_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16238__A3 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17862_ _17894_/A _17862_/B _17862_/C VGND VGND VPWR VPWR _17866_/B sky130_fd_sc_hd__and3_4
XFILLER_61_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19601_ _21913_/B _19596_/X _19600_/X _19596_/X VGND VGND VPWR VPWR _19601_/X sky130_fd_sc_hd__a2bb2o_4
X_16813_ _17053_/A VGND VGND VPWR VPWR _17067_/A sky130_fd_sc_hd__buf_2
XANTENNA__17986__A3 _16096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17793_ _17929_/A _17791_/X _17792_/X VGND VGND VPWR VPWR _17793_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_204_0_HCLK clkbuf_8_205_0_HCLK/A VGND VGND VPWR VPWR _24171_/CLK sky130_fd_sc_hd__clkbuf_1
X_19532_ _19530_/X _18025_/D _19531_/X VGND VGND VPWR VPWR _19533_/A sky130_fd_sc_hd__or3_4
X_16744_ _16740_/X _16744_/B _16742_/X _16743_/X VGND VGND VPWR VPWR _16745_/D sky130_fd_sc_hd__or4_4
X_13956_ _13937_/A VGND VGND VPWR VPWR _13956_/X sky130_fd_sc_hd__buf_2
XFILLER_98_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12907_ _12907_/A VGND VGND VPWR VPWR _12908_/B sky130_fd_sc_hd__inv_2
X_19463_ _19461_/Y _19458_/X _19462_/X _19458_/X VGND VGND VPWR VPWR _23328_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13887_ _13887_/A _13886_/X VGND VGND VPWR VPWR _13887_/X sky130_fd_sc_hd__or2_4
X_16675_ _13461_/C VGND VGND VPWR VPWR _20919_/A sky130_fd_sc_hd__inv_2
XANTENNA__15749__A2 _15740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18414_ _23839_/Q VGND VGND VPWR VPWR _18438_/A sky130_fd_sc_hd__inv_2
X_12838_ _22769_/A VGND VGND VPWR VPWR _12838_/Y sky130_fd_sc_hd__inv_2
X_15626_ _12575_/Y _15624_/X _15386_/X _15624_/X VGND VGND VPWR VPWR _24509_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24486__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19394_ _13030_/B VGND VGND VPWR VPWR _19394_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18345_ _23838_/Q VGND VGND VPWR VPWR _18472_/A sky130_fd_sc_hd__buf_2
XFILLER_61_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24415__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12769_ _12735_/X VGND VGND VPWR VPWR _12770_/B sky130_fd_sc_hd__inv_2
X_15557_ _15556_/X VGND VGND VPWR VPWR _15557_/Y sky130_fd_sc_hd__inv_2
XPHY_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14508_ _14501_/X _14505_/Y _14507_/Y VGND VGND VPWR VPWR _14508_/X sky130_fd_sc_hd__a21o_4
XANTENNA_clkbuf_2_1_0_HCLK_A clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15488_ _12088_/Y _15487_/X _15350_/X _15487_/X VGND VGND VPWR VPWR _24566_/D sky130_fd_sc_hd__a2bb2o_4
X_18276_ _18205_/A _18280_/B _18275_/Y VGND VGND VPWR VPWR _23864_/D sky130_fd_sc_hd__o21a_4
XFILLER_30_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17227_ _23896_/Q _17227_/B VGND VGND VPWR VPWR _17228_/A sky130_fd_sc_hd__and2_4
X_14439_ _14541_/D VGND VGND VPWR VPWR _19904_/D sky130_fd_sc_hd__buf_2
XANTENNA__19448__A _19448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15382__B1 _11604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21455__B1 _11961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11538__A3 _11536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17158_ _17157_/X VGND VGND VPWR VPWR _24031_/D sky130_fd_sc_hd__inv_2
X_16109_ _24331_/Q VGND VGND VPWR VPWR _22014_/A sky130_fd_sc_hd__inv_2
XANTENNA__15134__B1 _15126_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17089_ _17089_/A _17092_/B VGND VGND VPWR VPWR _17090_/C sky130_fd_sc_hd__or2_4
XFILLER_89_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11728__B _11720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22602__A _16172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_14_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_14_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__25203__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22321__B _22320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16634__B1 _22857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13448__B1 _13446_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22707__B1 _25211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22810_ _22810_/A _22884_/B VGND VGND VPWR VPWR _22810_/X sky130_fd_sc_hd__and2_4
X_23790_ _24811_/CLK _11916_/C HRESETn VGND VGND VPWR VPWR _11910_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_77_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22741_ _22539_/X _22739_/X _20750_/X _22740_/Y VGND VGND VPWR VPWR _22742_/A sky130_fd_sc_hd__o22a_4
XFILLER_37_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_1_HCLK clkbuf_1_0_1_HCLK/A VGND VGND VPWR VPWR clkbuf_2_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22672_ _22547_/X _22670_/X _22551_/X _22671_/X VGND VGND VPWR VPWR _22673_/B sky130_fd_sc_hd__o22a_4
XANTENNA__22049__A _21490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24411_ _24412_/CLK _15869_/X HRESETn VGND VGND VPWR VPWR _24411_/Q sky130_fd_sc_hd__dfrtp_4
X_21623_ _18043_/A _21621_/X _21622_/X VGND VGND VPWR VPWR _21623_/X sky130_fd_sc_hd__and3_4
XANTENNA__24156__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24342_ _23872_/CLK _24342_/D HRESETn VGND VGND VPWR VPWR _16078_/A sky130_fd_sc_hd__dfrtp_4
X_21554_ _21860_/B VGND VGND VPWR VPWR _22227_/B sky130_fd_sc_hd__buf_2
X_20505_ _22624_/A _20416_/A _20446_/X _20504_/Y VGND VGND VPWR VPWR _20506_/A sky130_fd_sc_hd__o22a_4
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24273_ _24676_/CLK _24273_/D HRESETn VGND VGND VPWR VPWR _24273_/Q sky130_fd_sc_hd__dfrtp_4
X_21485_ _21352_/A _19293_/Y VGND VGND VPWR VPWR _21485_/X sky130_fd_sc_hd__or2_4
XFILLER_5_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23224_ _23401_/CLK _19753_/X VGND VGND VPWR VPWR _19752_/A sky130_fd_sc_hd__dfxtp_4
X_20436_ _20436_/A VGND VGND VPWR VPWR _20436_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23155_ _23154_/CLK _23155_/D VGND VGND VPWR VPWR _23155_/Q sky130_fd_sc_hd__dfxtp_4
X_20367_ _20343_/Y VGND VGND VPWR VPWR _20367_/X sky130_fd_sc_hd__buf_2
XFILLER_101_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23791__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22106_ _20964_/A _22106_/B VGND VGND VPWR VPWR _22108_/B sky130_fd_sc_hd__or2_4
XANTENNA__23720__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23086_ _23383_/CLK _23086_/D VGND VGND VPWR VPWR _20114_/A sky130_fd_sc_hd__dfxtp_4
X_20298_ _20298_/A _20297_/Y _20278_/X VGND VGND VPWR VPWR _20298_/X sky130_fd_sc_hd__and3_4
XANTENNA__22512__A _22512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21749__A1 _13428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22946__B1 _13362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22037_ _14618_/A _22246_/B _14077_/A _21357_/A VGND VGND VPWR VPWR _22037_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17606__A _16685_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24997__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13810_ _13810_/A VGND VGND VPWR VPWR _13810_/X sky130_fd_sc_hd__buf_2
X_14790_ _24688_/Q VGND VGND VPWR VPWR _15078_/A sky130_fd_sc_hd__inv_2
XFILLER_60_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24926__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23988_ _23986_/CLK _23988_/D HRESETn VGND VGND VPWR VPWR _17244_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_113_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22174__B2 _22173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13741_ _13722_/X _24635_/Q _13737_/A _13718_/X VGND VGND VPWR VPWR _13742_/D sky130_fd_sc_hd__or4_4
XFILLER_44_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22939_ _22919_/X _22923_/X _22938_/X VGND VGND VPWR VPWR HRDATA[28] sky130_fd_sc_hd__a21o_4
XFILLER_113_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_34_0_HCLK clkbuf_8_35_0_HCLK/A VGND VGND VPWR VPWR _23401_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_5_18_0_HCLK_A clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13672_ _13419_/Y _13667_/X _13635_/X _13671_/X VGND VGND VPWR VPWR _24928_/D sky130_fd_sc_hd__a2bb2o_4
X_16460_ _16452_/A VGND VGND VPWR VPWR _16460_/X sky130_fd_sc_hd__buf_2
XFILLER_16_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_97_0_HCLK clkbuf_7_48_0_HCLK/X VGND VGND VPWR VPWR _24088_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12623_ _25040_/Q VGND VGND VPWR VPWR _12629_/A sky130_fd_sc_hd__inv_2
X_15411_ _15410_/X VGND VGND VPWR VPWR _15411_/X sky130_fd_sc_hd__buf_2
XFILLER_31_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16391_ _21109_/B VGND VGND VPWR VPWR _21047_/A sky130_fd_sc_hd__buf_2
XFILLER_58_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24609_ _24182_/CLK _24609_/D HRESETn VGND VGND VPWR VPWR _15339_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21449__A2_N _14015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15342_ _24608_/Q VGND VGND VPWR VPWR _15342_/Y sky130_fd_sc_hd__inv_2
X_18130_ _20736_/B VGND VGND VPWR VPWR _18130_/Y sky130_fd_sc_hd__inv_2
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12554_ _12553_/Y VGND VGND VPWR VPWR _12554_/X sky130_fd_sc_hd__buf_2
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11505_ _11505_/A VGND VGND VPWR VPWR _11507_/A sky130_fd_sc_hd__inv_2
XFILLER_78_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15273_ _15270_/Y _15272_/X _14228_/X _15272_/X VGND VGND VPWR VPWR _15273_/X sky130_fd_sc_hd__a2bb2o_4
X_18061_ _17446_/X _18061_/B _18060_/X VGND VGND VPWR VPWR _18061_/X sky130_fd_sc_hd__or3_4
XFILLER_89_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15364__B1 _11576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12485_ _12485_/A VGND VGND VPWR VPWR _12485_/Y sky130_fd_sc_hd__inv_2
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23879__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14224_ _14196_/X VGND VGND VPWR VPWR _18633_/A sky130_fd_sc_hd__buf_2
X_17012_ _17005_/X _17007_/X _17012_/C _17012_/D VGND VGND VPWR VPWR _17012_/X sky130_fd_sc_hd__or4_4
XFILLER_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21988__A1 _22155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14155_ _18111_/B _14153_/X VGND VGND VPWR VPWR _14155_/X sky130_fd_sc_hd__or2_4
XFILLER_98_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18900__A _18899_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13106_ _13309_/A _13106_/B VGND VGND VPWR VPWR _13106_/X sky130_fd_sc_hd__or2_4
XFILLER_3_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14086_ _24859_/Q VGND VGND VPWR VPWR _14086_/Y sky130_fd_sc_hd__inv_2
X_18963_ _18963_/A VGND VGND VPWR VPWR _18963_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13037_ _11735_/Y VGND VGND VPWR VPWR _13113_/A sky130_fd_sc_hd__buf_2
X_17914_ _17914_/A _17912_/X _17914_/C VGND VGND VPWR VPWR _17915_/C sky130_fd_sc_hd__and3_4
X_18894_ _18893_/Y _18891_/X _18802_/X _18891_/X VGND VGND VPWR VPWR _18894_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16420__A _24211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15419__A1 _15411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12350__B1 _12534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17845_ _17877_/A _17845_/B VGND VGND VPWR VPWR _17845_/X sky130_fd_sc_hd__or2_4
XFILLER_113_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12080__A2_N _24570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21980__B _21979_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24667__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17776_ _17716_/X _17774_/X _17776_/C VGND VGND VPWR VPWR _17777_/C sky130_fd_sc_hd__and3_4
XFILLER_54_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14988_ _14990_/B VGND VGND VPWR VPWR _14989_/B sky130_fd_sc_hd__inv_2
X_19515_ _23308_/Q VGND VGND VPWR VPWR _19515_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16727_ _15968_/Y _22395_/A _15968_/Y _22395_/A VGND VGND VPWR VPWR _16731_/A sky130_fd_sc_hd__a2bb2o_4
X_13939_ _13939_/A VGND VGND VPWR VPWR _13939_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20028__A2_N _20027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19446_ _21942_/B _19441_/X _19445_/X _19441_/X VGND VGND VPWR VPWR _19446_/X sky130_fd_sc_hd__a2bb2o_4
X_16658_ _16658_/A VGND VGND VPWR VPWR _16658_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15609_ _12588_/Y _15607_/X _11570_/X _15607_/X VGND VGND VPWR VPWR _15609_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_5_5_0_HCLK clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19377_ _13144_/B VGND VGND VPWR VPWR _19377_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16589_ _16581_/X _16573_/X HWDATA[19] _24144_/Q _16566_/X VGND VGND VPWR VPWR _16589_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_128_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18328_ _18300_/A _18327_/X VGND VGND VPWR VPWR _18328_/Y sky130_fd_sc_hd__nand2_4
X_18259_ _18219_/X _18258_/X _18240_/C VGND VGND VPWR VPWR _18259_/X sky130_fd_sc_hd__o21a_4
XFILLER_129_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21270_ _15322_/A _21269_/X _21058_/X _12585_/A _21059_/X VGND VGND VPWR VPWR _21270_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15370__A3 _15369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20221_ _20232_/A _20221_/B _20220_/Y VGND VGND VPWR VPWR _20221_/X sky130_fd_sc_hd__or3_4
XFILLER_104_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20152_ _23069_/Q VGND VGND VPWR VPWR _20152_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13669__B1 _13668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14330__A1 _20331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24960_ _24957_/CLK _24960_/D HRESETn VGND VGND VPWR VPWR _13566_/C sky130_fd_sc_hd__dfrtp_4
X_20083_ _20081_/Y _20077_/X _19603_/A _20082_/X VGND VGND VPWR VPWR _20083_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16607__B1 _16455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23911_ _24928_/CLK _23911_/D HRESETn VGND VGND VPWR VPWR _11677_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_135_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24891_ _24783_/CLK _24891_/D HRESETn VGND VGND VPWR VPWR _24891_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17280__B1 _25211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23842_ _23824_/CLK _23842_/D HRESETn VGND VGND VPWR VPWR _23842_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20787__A _24360_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24337__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_250_0_HCLK clkbuf_8_251_0_HCLK/A VGND VGND VPWR VPWR _24112_/CLK sky130_fd_sc_hd__clkbuf_1
X_23773_ _24643_/CLK _20233_/X HRESETn VGND VGND VPWR VPWR _23773_/Q sky130_fd_sc_hd__dfrtp_4
X_20985_ _20978_/A _19571_/Y _17644_/A VGND VGND VPWR VPWR _20985_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21903__B2 _21088_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22724_ _16418_/Y _22551_/A _14781_/Y _22225_/A VGND VGND VPWR VPWR _22724_/X sky130_fd_sc_hd__o22a_4
XFILLER_53_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12601__A2_N _24516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15594__B1 _11540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22655_ _23961_/Q _22654_/X _22608_/X VGND VGND VPWR VPWR _22655_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21606_ _18043_/A _21603_/X _21605_/X VGND VGND VPWR VPWR _21606_/X sky130_fd_sc_hd__and3_4
X_22586_ _16510_/Y _22435_/X VGND VGND VPWR VPWR _22586_/X sky130_fd_sc_hd__and2_4
X_24325_ _24013_/CLK _24325_/D HRESETn VGND VGND VPWR VPWR _16123_/A sky130_fd_sc_hd__dfrtp_4
X_21537_ _21530_/Y _21536_/Y _21793_/A VGND VGND VPWR VPWR _21537_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15346__B1 _11555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23972__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20890__A1 _20885_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25196__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12270_ _12097_/Y _12282_/B VGND VGND VPWR VPWR _12280_/B sky130_fd_sc_hd__or2_4
X_24256_ _24262_/CLK _16293_/X HRESETn VGND VGND VPWR VPWR _14936_/A sky130_fd_sc_hd__dfrtp_4
X_21468_ _21144_/A _21466_/X _21468_/C VGND VGND VPWR VPWR _21468_/X sky130_fd_sc_hd__and3_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23901__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25125__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23207_ _25112_/CLK _23207_/D VGND VGND VPWR VPWR _23207_/Q sky130_fd_sc_hd__dfxtp_4
X_20419_ _20511_/A VGND VGND VPWR VPWR _20419_/X sky130_fd_sc_hd__buf_2
X_24187_ _24185_/CLK _24187_/D HRESETn VGND VGND VPWR VPWR _24187_/Q sky130_fd_sc_hd__dfrtp_4
X_21399_ _20892_/X _21398_/X _13637_/A _22548_/A VGND VGND VPWR VPWR _21399_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15649__A1 _15411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23138_ _23313_/CLK _19980_/X VGND VGND VPWR VPWR _19979_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_134_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15960_ _15921_/X VGND VGND VPWR VPWR _15987_/A sky130_fd_sc_hd__buf_2
X_23069_ _23992_/CLK _23069_/D VGND VGND VPWR VPWR _23069_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_103_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14911_ _24658_/Q _24263_/Q _15108_/B _14910_/Y VGND VGND VPWR VPWR _14911_/X sky130_fd_sc_hd__o22a_4
X_15891_ _15889_/Y _15885_/X _15890_/X _15885_/X VGND VGND VPWR VPWR _15891_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_6_60_0_HCLK clkbuf_6_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_60_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17630_ _23940_/Q _17630_/B VGND VGND VPWR VPWR _17632_/A sky130_fd_sc_hd__and2_4
X_14842_ _15004_/A _24148_/Q _15004_/A _24148_/Q VGND VGND VPWR VPWR _14842_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24760__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14085__B1 _13668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17561_ _17498_/Y _17550_/B VGND VGND VPWR VPWR _17565_/A sky130_fd_sc_hd__or2_4
XFILLER_112_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24078__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11985_ _25147_/Q VGND VGND VPWR VPWR _11985_/Y sky130_fd_sc_hd__inv_2
X_14773_ _14764_/X _14773_/B _14769_/X _14772_/X VGND VGND VPWR VPWR _14794_/B sky130_fd_sc_hd__or4_4
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19300_ _19300_/A VGND VGND VPWR VPWR _19300_/Y sky130_fd_sc_hd__inv_2
X_16512_ _16510_/Y _16506_/X _16264_/X _16511_/X VGND VGND VPWR VPWR _16512_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17071__A _17052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13724_ _24635_/Q VGND VGND VPWR VPWR _13745_/B sky130_fd_sc_hd__buf_2
XANTENNA__24007__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17492_ _17484_/Y _17486_/X _17489_/X _17492_/D VGND VGND VPWR VPWR _17492_/X sky130_fd_sc_hd__or4_4
X_19231_ _19231_/A VGND VGND VPWR VPWR _19231_/Y sky130_fd_sc_hd__inv_2
X_16443_ _16443_/A VGND VGND VPWR VPWR _16443_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13655_ _13655_/A VGND VGND VPWR VPWR _13655_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13104__A _13182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _12605_/Y _24525_/Q _12605_/Y _24525_/Q VGND VGND VPWR VPWR _12606_/X sky130_fd_sc_hd__a2bb2o_4
X_19162_ _23432_/Q VGND VGND VPWR VPWR _19162_/Y sky130_fd_sc_hd__inv_2
X_13586_ _13550_/Y VGND VGND VPWR VPWR _13586_/X sky130_fd_sc_hd__buf_2
X_16374_ _16371_/Y _16372_/X _16373_/X _16372_/X VGND VGND VPWR VPWR _16374_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18113_ _18118_/A VGND VGND VPWR VPWR _18113_/X sky130_fd_sc_hd__buf_2
X_12537_ _12456_/X _12537_/B _12537_/C VGND VGND VPWR VPWR _12537_/X sky130_fd_sc_hd__and3_4
X_15325_ _15325_/A VGND VGND VPWR VPWR _15401_/A sky130_fd_sc_hd__inv_2
XFILLER_125_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21311__A2_N _11503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19093_ _19091_/Y _19092_/X _18959_/X _19092_/X VGND VGND VPWR VPWR _23457_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18044_ _18030_/A _18038_/A _18033_/X VGND VGND VPWR VPWR _18044_/X sky130_fd_sc_hd__a21o_4
X_12468_ _12468_/A VGND VGND VPWR VPWR _12469_/B sky130_fd_sc_hd__inv_2
X_15256_ _15240_/A VGND VGND VPWR VPWR _15256_/X sky130_fd_sc_hd__buf_2
XANTENNA__23642__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14207_ _20188_/A _14200_/X _13668_/X _14202_/X VGND VGND VPWR VPWR _14207_/X sky130_fd_sc_hd__a2bb2o_4
X_15187_ _15123_/A _15187_/B VGND VGND VPWR VPWR _15188_/B sky130_fd_sc_hd__or2_4
X_12399_ _12399_/A VGND VGND VPWR VPWR _12434_/A sky130_fd_sc_hd__buf_2
X_14138_ _14126_/A _14137_/X _13348_/A _14131_/X VGND VGND VPWR VPWR _24844_/D sky130_fd_sc_hd__o22a_4
XFILLER_113_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14767__A2_N _24116_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19995_ _23132_/Q VGND VGND VPWR VPWR _19995_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14069_ _13792_/C _14068_/X VGND VGND VPWR VPWR _15251_/A sky130_fd_sc_hd__or2_4
X_18946_ _18942_/Y _18945_/X _18901_/X _18945_/X VGND VGND VPWR VPWR _23510_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24848__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18877_ _18876_/Y VGND VGND VPWR VPWR _18877_/X sky130_fd_sc_hd__buf_2
XFILLER_66_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17828_ _17895_/A _17828_/B VGND VGND VPWR VPWR _17830_/B sky130_fd_sc_hd__or2_4
XFILLER_55_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14076__B1 sda_oen_o_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24430__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17759_ _14571_/X _23517_/Q VGND VGND VPWR VPWR _17759_/X sky130_fd_sc_hd__or2_4
XANTENNA__20149__B1 _19808_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12626__B2 _24532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20770_ _20750_/X _20754_/X _20769_/X VGND VGND VPWR VPWR _20770_/X sky130_fd_sc_hd__and3_4
XFILLER_74_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19429_ _19429_/A VGND VGND VPWR VPWR _19429_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_80_0_HCLK clkbuf_8_81_0_HCLK/A VGND VGND VPWR VPWR _23648_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22440_ _16089_/Y _22859_/A VGND VGND VPWR VPWR _22441_/C sky130_fd_sc_hd__or2_4
XANTENNA__15328__B1 _11522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22371_ _22369_/X _22370_/X _21986_/X _24407_/Q _21987_/X VGND VGND VPWR VPWR _22371_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22861__A2 _15919_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24110_ _24698_/CLK _24110_/D HRESETn VGND VGND VPWR VPWR _14751_/A sky130_fd_sc_hd__dfrtp_4
X_21322_ _21322_/A VGND VGND VPWR VPWR _21323_/D sky130_fd_sc_hd__inv_2
XFILLER_50_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_0_0_HCLK clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_2_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_25090_ _25090_/CLK _12473_/Y HRESETn VGND VGND VPWR VPWR _22678_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_129_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24041_ _24042_/CLK _17122_/Y HRESETn VGND VGND VPWR VPWR _24041_/Q sky130_fd_sc_hd__dfrtp_4
X_21253_ _11941_/X _21251_/X _21252_/X _13641_/Y _21720_/B VGND VGND VPWR VPWR _21253_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19636__A _19636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20204_ _23658_/Q VGND VGND VPWR VPWR _20204_/X sky130_fd_sc_hd__buf_2
XANTENNA__21821__B1 _20968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21184_ _21184_/A VGND VGND VPWR VPWR _21184_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20135_ _20134_/X VGND VGND VPWR VPWR _20141_/A sky130_fd_sc_hd__inv_2
XANTENNA__17156__A _17086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18578__A1_N _24249_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15500__B1 _24559_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24589__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22997__A _22997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20066_ _23104_/Q VGND VGND VPWR VPWR _20066_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24518__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24943_ _24944_/CLK _24943_/D HRESETn VGND VGND VPWR VPWR _13637_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19242__B2 _19239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_4_0_HCLK_A clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18450__C1 _18449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24874_ _23657_/CLK _14040_/X HRESETn VGND VGND VPWR VPWR _24874_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24171__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23825_ _23826_/CLK _23825_/D HRESETn VGND VGND VPWR VPWR _23825_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17005__B1 _16193_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24100__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11770_ _17448_/A VGND VGND VPWR VPWR _11809_/A sky130_fd_sc_hd__buf_2
XFILLER_92_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23756_ _24185_/CLK _23756_/D HRESETn VGND VGND VPWR VPWR _23756_/Q sky130_fd_sc_hd__dfrtp_4
X_20968_ _23940_/Q VGND VGND VPWR VPWR _20968_/X sky130_fd_sc_hd__buf_2
XFILLER_92_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17556__A1 _17497_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22707_ _22369_/X _22706_/X _22640_/X _25211_/Q _22641_/X VGND VGND VPWR VPWR _22707_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20560__B1 _20556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23687_ _24879_/CLK _23687_/D HRESETn VGND VGND VPWR VPWR _23687_/Q sky130_fd_sc_hd__dfrtp_4
X_20899_ _21109_/B VGND VGND VPWR VPWR _20900_/A sky130_fd_sc_hd__buf_2
X_13440_ _13430_/X _13440_/B _13436_/X _13440_/D VGND VGND VPWR VPWR _13440_/X sky130_fd_sc_hd__or4_4
Xclkbuf_8_108_0_HCLK clkbuf_7_54_0_HCLK/X VGND VGND VPWR VPWR _24587_/CLK sky130_fd_sc_hd__clkbuf_1
X_22638_ _21293_/B VGND VGND VPWR VPWR _22638_/X sky130_fd_sc_hd__buf_2
XFILLER_16_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12555__A2_N _24518_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22237__A _21642_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22301__B2 _20866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13371_ _13370_/Y _13366_/X _11620_/X _13366_/X VGND VGND VPWR VPWR _24982_/D sky130_fd_sc_hd__a2bb2o_4
X_22569_ _20630_/Y _22279_/X _20495_/C _22322_/A VGND VGND VPWR VPWR _22569_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16235__A _22477_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12322_ _12322_/A VGND VGND VPWR VPWR _12405_/D sky130_fd_sc_hd__inv_2
X_15110_ _15224_/A _15110_/B _14883_/Y _15109_/Y VGND VGND VPWR VPWR _15110_/X sky130_fd_sc_hd__or4_4
XFILLER_126_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16090_ _16084_/A VGND VGND VPWR VPWR _16090_/X sky130_fd_sc_hd__buf_2
X_24308_ _24308_/CLK _16171_/X HRESETn VGND VGND VPWR VPWR _24308_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20980__A _20980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15041_ _15041_/A VGND VGND VPWR VPWR _24698_/D sky130_fd_sc_hd__inv_2
X_12253_ _12237_/A _12228_/X _12203_/X _12250_/Y VGND VGND VPWR VPWR _12254_/A sky130_fd_sc_hd__a211o_4
X_24239_ _23830_/CLK _16344_/X HRESETn VGND VGND VPWR VPWR _24239_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12184_ _12079_/X _12219_/A _12171_/X _12184_/D VGND VGND VPWR VPWR _12184_/X sky130_fd_sc_hd__or4_4
XFILLER_29_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18800_ _18800_/A VGND VGND VPWR VPWR _18800_/Y sky130_fd_sc_hd__inv_2
X_19780_ _19780_/A VGND VGND VPWR VPWR _19780_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24941__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16992_ _16992_/A VGND VGND VPWR VPWR _16992_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18731_ _18730_/Y _18719_/A _18712_/X _18719_/A VGND VGND VPWR VPWR _18731_/X sky130_fd_sc_hd__a2bb2o_4
X_15943_ _22763_/A VGND VGND VPWR VPWR _15943_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24259__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18662_ _19859_/A VGND VGND VPWR VPWR _18662_/X sky130_fd_sc_hd__buf_2
X_15874_ _15872_/Y _15868_/X _11585_/X _15873_/X VGND VGND VPWR VPWR _24409_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14058__B1 _13635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17613_ _17488_/Y _17510_/B VGND VGND VPWR VPWR _17614_/B sky130_fd_sc_hd__or2_4
X_14825_ _24155_/Q VGND VGND VPWR VPWR _14825_/Y sky130_fd_sc_hd__inv_2
X_18593_ _16371_/A _18543_/A _16358_/Y _18338_/X VGND VGND VPWR VPWR _18593_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12938__A _22712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17544_ _17502_/D _17511_/B _17502_/B VGND VGND VPWR VPWR _17544_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21879__B1 _13337_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14756_ _24683_/Q _14754_/Y _24687_/Q _14755_/Y VGND VGND VPWR VPWR _14761_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11968_ _25154_/Q VGND VGND VPWR VPWR _11968_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22540__A1 _12592_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22540__B2 _22029_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13707_ _13697_/X _13706_/X _24856_/Q _13682_/Y VGND VGND VPWR VPWR _24915_/D sky130_fd_sc_hd__o22a_4
X_17475_ _17474_/Y _17462_/Y _21801_/A _17461_/X VGND VGND VPWR VPWR _17475_/X sky130_fd_sc_hd__o22a_4
X_11899_ _11883_/A _11894_/A _11898_/Y VGND VGND VPWR VPWR _11900_/A sky130_fd_sc_hd__o21a_4
X_14687_ _14683_/A _14682_/X _14683_/Y VGND VGND VPWR VPWR _14687_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__23894__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_67_0_HCLK clkbuf_7_67_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_67_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19214_ _19211_/Y _19213_/X _19170_/X _19213_/X VGND VGND VPWR VPWR _19214_/X sky130_fd_sc_hd__a2bb2o_4
X_16426_ _16426_/A VGND VGND VPWR VPWR _16426_/X sky130_fd_sc_hd__buf_2
XFILLER_38_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13638_ _15801_/A VGND VGND VPWR VPWR _13638_/X sky130_fd_sc_hd__buf_2
XFILLER_20_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23823__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22147__A _22147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21051__A _21050_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25047__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19145_ _19144_/X VGND VGND VPWR VPWR _19153_/A sky130_fd_sc_hd__inv_2
X_16357_ _16356_/Y _16352_/X _16096_/X _16352_/X VGND VGND VPWR VPWR _16357_/X sky130_fd_sc_hd__a2bb2o_4
X_13569_ _13568_/X VGND VGND VPWR VPWR _13569_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16145__A _16165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12792__B1 _22900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15308_ _14013_/A VGND VGND VPWR VPWR _21300_/A sky130_fd_sc_hd__buf_2
X_19076_ _19075_/Y _19071_/X _18964_/X _19071_/A VGND VGND VPWR VPWR _23463_/D sky130_fd_sc_hd__a2bb2o_4
X_16288_ _15915_/X _16276_/X _15704_/X _24259_/Q _16237_/A VGND VGND VPWR VPWR _24259_/D
+ sky130_fd_sc_hd__a32o_4
X_18027_ _18023_/A VGND VGND VPWR VPWR _18031_/B sky130_fd_sc_hd__inv_2
XANTENNA__15984__A _24367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15239_ _15241_/A VGND VGND VPWR VPWR _15240_/A sky130_fd_sc_hd__buf_2
XFILLER_132_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19978_ _19977_/Y _19975_/X _19452_/A _19975_/X VGND VGND VPWR VPWR _19978_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24682__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22359__B2 _22358_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18929_ _17838_/B VGND VGND VPWR VPWR _18929_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12003__A1_N _12001_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24611__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22610__A _22610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_HCLK HCLK VGND VGND VPWR VPWR clkbuf_0_HCLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_67_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21940_ _21229_/A _21940_/B VGND VGND VPWR VPWR _21940_/X sky130_fd_sc_hd__or2_4
XFILLER_55_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14049__B1 _13663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18983__B1 _18959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21871_ _21871_/A _20885_/X VGND VGND VPWR VPWR _21871_/X sky130_fd_sc_hd__or2_4
XFILLER_54_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11752__A _11751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23610_ _23489_/CLK _18655_/X VGND VGND VPWR VPWR _18654_/A sky130_fd_sc_hd__dfxtp_4
X_20822_ _20822_/A _20821_/X VGND VGND VPWR VPWR _20822_/Y sky130_fd_sc_hd__nand2_4
XPHY_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24590_ _24590_/CLK _15391_/X HRESETn VGND VGND VPWR VPWR _24590_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23541_ _23133_/CLK _18857_/X VGND VGND VPWR VPWR _13063_/B sky130_fd_sc_hd__dfxtp_4
X_20753_ _20753_/A VGND VGND VPWR VPWR _23025_/B sky130_fd_sc_hd__buf_2
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23472_ _24998_/CLK _23472_/D VGND VGND VPWR VPWR _19051_/A sky130_fd_sc_hd__dfxtp_4
X_20684_ _24996_/Q _11706_/A _11708_/B VGND VGND VPWR VPWR _23781_/D sky130_fd_sc_hd__a21o_4
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25211_ _24590_/CLK _11561_/X HRESETn VGND VGND VPWR VPWR _25211_/Q sky130_fd_sc_hd__dfrtp_4
X_22423_ _21569_/A VGND VGND VPWR VPWR _22423_/X sky130_fd_sc_hd__buf_2
XANTENNA__21098__B2 _20863_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22295__B1 _25201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25142_ _23789_/CLK _25142_/D HRESETn VGND VGND VPWR VPWR _12001_/A sky130_fd_sc_hd__dfrtp_4
X_22354_ _22354_/A VGND VGND VPWR VPWR _22354_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21896__A _22228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21305_ _13326_/A _21303_/X _11954_/A _21304_/X VGND VGND VPWR VPWR _21305_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15894__A _16373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25073_ _25091_/CLK _25073_/D HRESETn VGND VGND VPWR VPWR _25073_/Q sky130_fd_sc_hd__dfrtp_4
X_22285_ _21020_/B VGND VGND VPWR VPWR _22285_/X sky130_fd_sc_hd__buf_2
XFILLER_3_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24024_ _23664_/CLK _24024_/D HRESETn VGND VGND VPWR VPWR _24024_/Q sky130_fd_sc_hd__dfstp_4
X_21236_ _21387_/A _21233_/X _21235_/X VGND VGND VPWR VPWR _21236_/X sky130_fd_sc_hd__and3_4
XANTENNA__16277__A1 _15915_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21270__A1 _15322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21167_ _21350_/A _21167_/B _21166_/X VGND VGND VPWR VPWR _21167_/X sky130_fd_sc_hd__and3_4
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14303__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20118_ _20054_/X _15641_/X _13663_/A _23085_/Q _20117_/X VGND VGND VPWR VPWR _20118_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24352__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21098_ _21719_/A _21097_/X _16385_/Y _20863_/A VGND VGND VPWR VPWR _21098_/X sky130_fd_sc_hd__o22a_4
XFILLER_58_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12940_ _12952_/A _12938_/X _12939_/X VGND VGND VPWR VPWR _12940_/X sky130_fd_sc_hd__and3_4
X_20049_ _21342_/B _20048_/X _19728_/X _20048_/X VGND VGND VPWR VPWR _20049_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17614__A _17614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24926_ _24928_/CLK _24926_/D HRESETn VGND VGND VPWR VPWR _24926_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21136__A _17651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12871_ _12781_/Y _12802_/Y VGND VGND VPWR VPWR _12884_/C sky130_fd_sc_hd__or2_4
X_24857_ _23657_/CLK _24857_/D HRESETn VGND VGND VPWR VPWR _14090_/A sky130_fd_sc_hd__dfrtp_4
X_14610_ _24719_/Q _14610_/B _14625_/A VGND VGND VPWR VPWR _14610_/X sky130_fd_sc_hd__or3_4
XFILLER_27_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11822_ _25178_/Q _11824_/A _11814_/Y _11821_/Y VGND VGND VPWR VPWR _11822_/X sky130_fd_sc_hd__o22a_4
X_23808_ _23648_/CLK _18628_/X HRESETn VGND VGND VPWR VPWR _23808_/Q sky130_fd_sc_hd__dfstp_4
X_15590_ _15593_/A VGND VGND VPWR VPWR _15590_/X sky130_fd_sc_hd__buf_2
XFILLER_45_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22522__A1 _22369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20975__A _20975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24788_ _24788_/CLK _14296_/X HRESETn VGND VGND VPWR VPWR _24788_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _11753_/A VGND VGND VPWR VPWR _13050_/A sky130_fd_sc_hd__buf_2
X_14541_ _14452_/X _14437_/X _14548_/A _14541_/D VGND VGND VPWR VPWR _14541_/X sky130_fd_sc_hd__and4_4
XFILLER_42_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20533__B1 _24610_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23739_ _24259_/CLK _20613_/X HRESETn VGND VGND VPWR VPWR _20611_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18445__A _18468_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _24007_/Q VGND VGND VPWR VPWR _17260_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _11683_/Y _23910_/Q _11683_/Y _23910_/Q VGND VGND VPWR VPWR _11693_/A sky130_fd_sc_hd__a2bb2o_4
X_14472_ _14469_/X VGND VGND VPWR VPWR _21396_/A sky130_fd_sc_hd__buf_2
XFILLER_41_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ _15282_/A VGND VGND VPWR VPWR _16211_/X sky130_fd_sc_hd__buf_2
XANTENNA__25140__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ _24762_/Q VGND VGND VPWR VPWR _14383_/A sky130_fd_sc_hd__inv_2
XANTENNA__21089__B2 _21088_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17191_ _17171_/X _17185_/X _23684_/Q _24024_/Q _17188_/X VGND VGND VPWR VPWR _24024_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14799__A1_N _15045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13354_ _13353_/Y _13351_/X _11981_/X _13351_/X VGND VGND VPWR VPWR _24988_/D sky130_fd_sc_hd__a2bb2o_4
X_16142_ _16140_/Y _16138_/X _16141_/X _16138_/X VGND VGND VPWR VPWR _24319_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12305_ _25101_/Q VGND VGND VPWR VPWR _12305_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13285_ _13221_/A _13283_/X _13284_/X VGND VGND VPWR VPWR _13285_/X sky130_fd_sc_hd__and3_4
X_16073_ _24344_/Q VGND VGND VPWR VPWR _16073_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12236_ _12235_/X VGND VGND VPWR VPWR _12236_/Y sky130_fd_sc_hd__inv_2
X_15024_ _14712_/X _15023_/Y VGND VGND VPWR VPWR _15024_/X sky130_fd_sc_hd__or2_4
X_19901_ _19901_/A VGND VGND VPWR VPWR _19901_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_9_0_HCLK clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19832_ _24536_/Q VGND VGND VPWR VPWR _19832_/X sky130_fd_sc_hd__buf_2
XANTENNA__21261__A1 _21247_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12167_ _24500_/Q VGND VGND VPWR VPWR _12167_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15309__A _21300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14213__A _15801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19763_ _19762_/Y _19760_/X _19714_/X _19760_/X VGND VGND VPWR VPWR _23221_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24093__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12098_ _12098_/A VGND VGND VPWR VPWR _12098_/Y sky130_fd_sc_hd__inv_2
X_16975_ _22164_/A VGND VGND VPWR VPWR _17145_/A sky130_fd_sc_hd__inv_2
XANTENNA__22430__A _15655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13474__D _21257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18714_ _17701_/B VGND VGND VPWR VPWR _18714_/Y sky130_fd_sc_hd__inv_2
X_15926_ _15925_/Y _15923_/X _11522_/X _15923_/X VGND VGND VPWR VPWR _15926_/X sky130_fd_sc_hd__a2bb2o_4
X_19694_ _19688_/Y VGND VGND VPWR VPWR _19694_/X sky130_fd_sc_hd__buf_2
XANTENNA__18965__B1 _18964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_30_0_HCLK clkbuf_5_30_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_61_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__22761__B2 _21187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18645_ _18644_/Y VGND VGND VPWR VPWR _18645_/X sky130_fd_sc_hd__buf_2
X_15857_ _24415_/Q VGND VGND VPWR VPWR _15857_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11572__A _25207_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14808_ _14791_/X _24128_/Q _14791_/X _24128_/Q VGND VGND VPWR VPWR _14808_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18576_ _18576_/A _18573_/X _18574_/X _18575_/X VGND VGND VPWR VPWR _18576_/X sky130_fd_sc_hd__or4_4
X_15788_ _15788_/A VGND VGND VPWR VPWR _15788_/X sky130_fd_sc_hd__buf_2
XFILLER_91_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18717__B1 _17202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17527_ _17509_/A _17525_/X _17526_/X VGND VGND VPWR VPWR _17527_/X sky130_fd_sc_hd__and3_4
X_14739_ _24711_/Q VGND VGND VPWR VPWR _14990_/A sky130_fd_sc_hd__inv_2
XFILLER_32_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19390__B1 _19366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17458_ _17455_/Y _17453_/X _17457_/Y VGND VGND VPWR VPWR _17458_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__14203__B1 _13663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16409_ _16426_/A VGND VGND VPWR VPWR _16409_/X sky130_fd_sc_hd__buf_2
X_17389_ _17270_/Y _17386_/B VGND VGND VPWR VPWR _17389_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15951__B1 _15770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19128_ _19127_/Y _19125_/X _19038_/X _19125_/X VGND VGND VPWR VPWR _23445_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_154_0_HCLK clkbuf_7_77_0_HCLK/X VGND VGND VPWR VPWR _25046_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_9_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19059_ _18763_/X VGND VGND VPWR VPWR _19059_/X sky130_fd_sc_hd__buf_2
XANTENNA__15703__B1 _15393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22324__B _22488_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22070_ _21665_/A _22068_/X _22070_/C VGND VGND VPWR VPWR _22074_/B sky130_fd_sc_hd__and3_4
XFILLER_82_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21021_ _15413_/A VGND VGND VPWR VPWR _21069_/A sky130_fd_sc_hd__inv_2
XFILLER_0_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22972_ _24459_/Q _22015_/X VGND VGND VPWR VPWR _22972_/X sky130_fd_sc_hd__or2_4
XFILLER_67_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18956__B1 _18932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24711_ _24671_/CLK _14991_/X HRESETn VGND VGND VPWR VPWR _24711_/Q sky130_fd_sc_hd__dfrtp_4
X_21923_ _17636_/X _21915_/X _21922_/X VGND VGND VPWR VPWR _21923_/X sky130_fd_sc_hd__and3_4
XFILLER_16_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21854_ _21051_/X _21853_/X VGND VGND VPWR VPWR _21855_/D sky130_fd_sc_hd__and2_4
X_24642_ _24644_/CLK _15258_/X HRESETn VGND VGND VPWR VPWR _13716_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_35_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23745__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15785__A3 _15505_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20805_ _20802_/X _20804_/X _12540_/Y _20802_/X VGND VGND VPWR VPWR _20805_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_70_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15889__A _15889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21785_ _21009_/A VGND VGND VPWR VPWR _21786_/A sky130_fd_sc_hd__buf_2
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24573_ _24573_/CLK _15474_/X HRESETn VGND VGND VPWR VPWR _24573_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20736_ _20736_/A _20736_/B VGND VGND VPWR VPWR _20736_/X sky130_fd_sc_hd__and2_4
XFILLER_24_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23524_ _23531_/CLK _18907_/X VGND VGND VPWR VPWR _23524_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_50_0_HCLK clkbuf_7_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_50_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22218__C _22218_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13548__A2 _20881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23455_ _23568_/CLK _23455_/D VGND VGND VPWR VPWR _23455_/Q sky130_fd_sc_hd__dfxtp_4
X_20667_ _23753_/Q _20664_/X _13539_/X VGND VGND VPWR VPWR _20667_/Y sky130_fd_sc_hd__a21boi_4
XANTENNA__15942__B1 _15761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19133__B1 _19109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22406_ _16559_/A _22405_/X VGND VGND VPWR VPWR _22416_/B sky130_fd_sc_hd__nor2_4
XFILLER_52_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23386_ _23112_/CLK _23386_/D VGND VGND VPWR VPWR _23386_/Q sky130_fd_sc_hd__dfxtp_4
X_20598_ _20647_/A VGND VGND VPWR VPWR _20598_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22337_ _21276_/A VGND VGND VPWR VPWR _22338_/A sky130_fd_sc_hd__buf_2
X_25125_ _25130_/CLK _12223_/X HRESETn VGND VGND VPWR VPWR _25125_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17609__A _23947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13070_ _13169_/A VGND VGND VPWR VPWR _13230_/A sky130_fd_sc_hd__buf_2
X_25056_ _24521_/CLK _25056_/D HRESETn VGND VGND VPWR VPWR _25056_/Q sky130_fd_sc_hd__dfrtp_4
X_22268_ _22264_/X _22267_/X _16361_/Y _13619_/X VGND VGND VPWR VPWR _22268_/X sky130_fd_sc_hd__o22a_4
XFILLER_2_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24533__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12021_ _12013_/A _23794_/Q _12020_/Y VGND VGND VPWR VPWR _12022_/A sky130_fd_sc_hd__o21a_4
XFILLER_65_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21725__A2_N _11954_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24007_ _24005_/CLK _17344_/X HRESETn VGND VGND VPWR VPWR _24007_/Q sky130_fd_sc_hd__dfrtp_4
X_21219_ _21237_/A VGND VGND VPWR VPWR _21224_/A sky130_fd_sc_hd__buf_2
X_22199_ _22195_/X _22196_/X _22197_/X _24404_/Q _22198_/X VGND VGND VPWR VPWR _22199_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_78_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22991__B2 _21561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22250__A _24477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16760_ _16760_/A VGND VGND VPWR VPWR _16760_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13972_ _13952_/X _13970_/Y _24890_/Q _13971_/X VGND VGND VPWR VPWR _13972_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15711_ _15693_/X _15460_/X _15635_/X _20808_/A _15661_/A VGND VGND VPWR VPWR _15711_/X
+ sky130_fd_sc_hd__a32o_4
X_12923_ _12802_/Y _12917_/B _12922_/X _12919_/B VGND VGND VPWR VPWR _12923_/X sky130_fd_sc_hd__a211o_4
XFILLER_47_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24909_ _24904_/CLK _24909_/D HRESETn VGND VGND VPWR VPWR _13828_/A sky130_fd_sc_hd__dfrtp_4
X_16691_ _22239_/A _17490_/A _15935_/Y _22853_/A VGND VGND VPWR VPWR _16691_/X sky130_fd_sc_hd__a2bb2o_4
X_18430_ _18430_/A VGND VGND VPWR VPWR _18430_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15642_ _15637_/X VGND VGND VPWR VPWR _15642_/X sky130_fd_sc_hd__buf_2
X_12854_ _12854_/A VGND VGND VPWR VPWR _12854_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11805_ _25180_/Q _11777_/X _13551_/B _11804_/Y VGND VGND VPWR VPWR _11805_/X sky130_fd_sc_hd__and4_4
X_18361_ _18361_/A VGND VGND VPWR VPWR _18536_/A sky130_fd_sc_hd__buf_2
XANTENNA__15799__A _16581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15573_ _22223_/A VGND VGND VPWR VPWR _16624_/A sky130_fd_sc_hd__buf_2
X_12785_ _12785_/A VGND VGND VPWR VPWR _12943_/C sky130_fd_sc_hd__buf_2
XPHY_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _17251_/Y _17382_/C _17312_/C _17311_/Y VGND VGND VPWR VPWR _17312_/X sky130_fd_sc_hd__or4_4
XANTENNA__22409__B _22488_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14524_ _14524_/A _14524_/B _14521_/X _14524_/D VGND VGND VPWR VPWR _14524_/X sky130_fd_sc_hd__and4_4
XFILLER_15_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11736_ _23897_/Q _23893_/Q _11734_/Y _11735_/Y VGND VGND VPWR VPWR _11738_/A sky130_fd_sc_hd__o22a_4
X_18292_ _18218_/B _18292_/B VGND VGND VPWR VPWR _18295_/B sky130_fd_sc_hd__or2_4
XPHY_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15528__A3 _15432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _11575_/Y _17309_/A _11575_/Y _17309_/A VGND VGND VPWR VPWR _17250_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ _21010_/A VGND VGND VPWR VPWR _21237_/A sky130_fd_sc_hd__buf_2
XFILLER_35_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11667_ _13566_/D VGND VGND VPWR VPWR _11667_/Y sky130_fd_sc_hd__inv_2
XPHY_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20809__A1 _20757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _13406_/A _13406_/B _13406_/C VGND VGND VPWR VPWR _13407_/B sky130_fd_sc_hd__and3_4
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17174_ _17174_/A _17174_/B VGND VGND VPWR VPWR _17174_/X sky130_fd_sc_hd__or2_4
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11598_ _16100_/A VGND VGND VPWR VPWR _11598_/X sky130_fd_sc_hd__buf_2
X_14386_ _14386_/A VGND VGND VPWR VPWR _14386_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15030__C _15033_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_227_0_HCLK clkbuf_8_227_0_HCLK/A VGND VGND VPWR VPWR _24308_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_127_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16125_ _24324_/Q VGND VGND VPWR VPWR _16125_/Y sky130_fd_sc_hd__inv_2
X_13337_ _13337_/A VGND VGND VPWR VPWR _14047_/A sky130_fd_sc_hd__buf_2
XFILLER_6_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_7_0_HCLK_A clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12951__A _12951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16056_ _16056_/A VGND VGND VPWR VPWR _16056_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24274__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13268_ _13300_/A _18684_/A VGND VGND VPWR VPWR _13270_/B sky130_fd_sc_hd__or2_4
XFILLER_131_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15007_ _24707_/Q _15006_/Y VGND VGND VPWR VPWR _15009_/B sky130_fd_sc_hd__or2_4
XFILLER_29_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12219_ _12219_/A _12219_/B VGND VGND VPWR VPWR _12219_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24203__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13199_ _13159_/X _13197_/X _13198_/X VGND VGND VPWR VPWR _13200_/C sky130_fd_sc_hd__and3_4
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19815_ _24541_/Q VGND VGND VPWR VPWR _19815_/X sky130_fd_sc_hd__buf_2
XANTENNA__16110__B1 _15890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16687__A2_N _17482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16958_ _16958_/A VGND VGND VPWR VPWR _24059_/D sky130_fd_sc_hd__inv_2
X_19746_ _21629_/B _19743_/X _19721_/X _19743_/X VGND VGND VPWR VPWR _23227_/D sky130_fd_sc_hd__a2bb2o_4
X_15909_ _15908_/Y _15826_/X _15291_/X _15826_/X VGND VGND VPWR VPWR _15909_/X sky130_fd_sc_hd__a2bb2o_4
X_19677_ _19677_/A VGND VGND VPWR VPWR _19677_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16889_ _16760_/Y _16887_/A VGND VGND VPWR VPWR _16889_/X sky130_fd_sc_hd__or2_4
XFILLER_65_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18628_ _18607_/X _18621_/X _23807_/Q _23808_/Q _18624_/X VGND VGND VPWR VPWR _18628_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25062__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18559_ _18355_/X _18559_/B VGND VGND VPWR VPWR _18559_/X sky130_fd_sc_hd__or2_4
XFILLER_21_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22319__B _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21570_ _21570_/A VGND VGND VPWR VPWR _21570_/X sky130_fd_sc_hd__buf_2
XFILLER_33_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_37_0_HCLK clkbuf_6_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_74_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20521_ _20520_/Y _20517_/Y _20524_/B VGND VGND VPWR VPWR _20521_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15924__B1 _15828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23240_ _23385_/CLK _19704_/X VGND VGND VPWR VPWR _23240_/Q sky130_fd_sc_hd__dfxtp_4
X_20452_ _20451_/X VGND VGND VPWR VPWR _23702_/D sky130_fd_sc_hd__inv_2
XFILLER_88_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22335__A _22335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23171_ _23156_/CLK _23171_/D VGND VGND VPWR VPWR _23171_/Q sky130_fd_sc_hd__dfxtp_4
X_20383_ _15284_/Y _20367_/X _20357_/X _20382_/X VGND VGND VPWR VPWR _20383_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22670__B1 _14958_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16333__A _16339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22122_ _22121_/X VGND VGND VPWR VPWR _22677_/A sky130_fd_sc_hd__buf_2
XFILLER_134_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22053_ _22064_/A _22053_/B VGND VGND VPWR VPWR _22053_/X sky130_fd_sc_hd__or2_4
XFILLER_121_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21004_ _21000_/X _21003_/X _24745_/Q VGND VGND VPWR VPWR _21004_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_134_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22973__A1 _23026_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22973__B2 _22460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16101__B1 _16100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23997__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22725__A1 _21529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23926__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22725__B2 _22724_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22955_ _22167_/A _22955_/B _22955_/C VGND VGND VPWR VPWR _22955_/X sky130_fd_sc_hd__and3_4
XFILLER_16_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21906_ _22806_/B _21896_/X _21900_/Y _21080_/Y _21905_/X VGND VGND VPWR VPWR _21906_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_55_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_119_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_239_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22886_ _22885_/X VGND VGND VPWR VPWR _22886_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21414__A _24432_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24625_ _24870_/CLK _15292_/X HRESETn VGND VGND VPWR VPWR _15290_/A sky130_fd_sc_hd__dfstp_4
X_21837_ _20750_/X _21798_/X _21807_/Y _20782_/X _21836_/X VGND VGND VPWR VPWR _21837_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12570_ _12568_/A _24510_/Q _12647_/B _12569_/Y VGND VGND VPWR VPWR _12570_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21768_ _21764_/X _21767_/X _14487_/X VGND VGND VPWR VPWR _21768_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__16168__B1 _15770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24556_ _25084_/CLK _15508_/X HRESETn VGND VGND VPWR VPWR _24556_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ _11521_/A VGND VGND VPWR VPWR _11521_/X sky130_fd_sc_hd__buf_2
X_20719_ _20719_/A _14023_/X VGND VGND VPWR VPWR _20719_/X sky130_fd_sc_hd__and2_4
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23507_ _23514_/CLK _23507_/D VGND VGND VPWR VPWR _17839_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_71_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14718__B2 _24093_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24785__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21699_ _21700_/A _21756_/B _13403_/Y _23393_/Q VGND VGND VPWR VPWR _21699_/X sky130_fd_sc_hd__o22a_4
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24487_ _25090_/CLK _24487_/D HRESETn VGND VGND VPWR VPWR _12382_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12474__C _12474_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14240_ _14239_/Y _14237_/X _14209_/X _14237_/X VGND VGND VPWR VPWR _14240_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24714__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23438_ _24735_/CLK _19147_/X VGND VGND VPWR VPWR _17697_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14171_ _14169_/B VGND VGND VPWR VPWR _14171_/X sky130_fd_sc_hd__buf_2
X_23369_ _24998_/CLK _23369_/D VGND VGND VPWR VPWR _13241_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA_clkbuf_5_0_0_HCLK_A clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16243__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13122_ _13122_/A _13119_/X _13121_/X VGND VGND VPWR VPWR _13122_/X sky130_fd_sc_hd__and3_4
X_25108_ _25115_/CLK _12285_/X HRESETn VGND VGND VPWR VPWR _25108_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16340__B1 _16261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_57_0_HCLK clkbuf_7_28_0_HCLK/X VGND VGND VPWR VPWR _24005_/CLK sky130_fd_sc_hd__clkbuf_1
X_13053_ _13053_/A _11648_/X _13053_/C VGND VGND VPWR VPWR _13053_/X sky130_fd_sc_hd__and3_4
X_17930_ _17815_/A _17930_/B _17929_/X VGND VGND VPWR VPWR _17938_/B sky130_fd_sc_hd__or3_4
XFILLER_79_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22413__B1 _16655_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25039_ _25009_/CLK _12768_/X HRESETn VGND VGND VPWR VPWR _12584_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23808__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12004_ _12004_/A VGND VGND VPWR VPWR _12004_/Y sky130_fd_sc_hd__inv_2
X_17861_ _17861_/A _17861_/B VGND VGND VPWR VPWR _17862_/C sky130_fd_sc_hd__or2_4
XFILLER_26_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16812_ _17132_/A VGND VGND VPWR VPWR _17053_/A sky130_fd_sc_hd__buf_2
X_19600_ _19600_/A VGND VGND VPWR VPWR _19600_/X sky130_fd_sc_hd__buf_2
XFILLER_78_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17792_ _17935_/A _18742_/A VGND VGND VPWR VPWR _17792_/X sky130_fd_sc_hd__or2_4
XFILLER_120_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23667__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19531_ _19531_/A _18022_/A _17625_/A VGND VGND VPWR VPWR _19531_/X sky130_fd_sc_hd__or3_4
X_16743_ _15986_/Y _16685_/A _15995_/Y _23945_/Q VGND VGND VPWR VPWR _16743_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13955_ _24806_/Q VGND VGND VPWR VPWR _13955_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12906_ _12963_/A _12885_/X VGND VGND VPWR VPWR _12907_/A sky130_fd_sc_hd__or2_4
X_19462_ _15561_/X VGND VGND VPWR VPWR _19462_/X sky130_fd_sc_hd__buf_2
XANTENNA__17802__A _16678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13107__A _13102_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16674_ _16652_/X _16653_/X _16558_/X _24093_/Q _16627_/A VGND VGND VPWR VPWR _24093_/D
+ sky130_fd_sc_hd__a32o_4
X_13886_ _13886_/A VGND VGND VPWR VPWR _13886_/X sky130_fd_sc_hd__buf_2
XFILLER_61_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15749__A3 _15468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18413_ _18413_/A VGND VGND VPWR VPWR _18462_/A sky130_fd_sc_hd__buf_2
X_15625_ _12569_/Y _15621_/X _15513_/X _15624_/X VGND VGND VPWR VPWR _15625_/X sky130_fd_sc_hd__a2bb2o_4
X_12837_ _12836_/Y _22385_/A _12836_/Y _22385_/A VGND VGND VPWR VPWR _12837_/X sky130_fd_sc_hd__a2bb2o_4
X_19393_ _19391_/Y _19386_/X _19392_/X _19372_/Y VGND VGND VPWR VPWR _23351_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18344_ _24196_/Q _18543_/A _16406_/Y _23840_/Q VGND VGND VPWR VPWR _18344_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15322__A _15322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15556_ _24536_/Q VGND VGND VPWR VPWR _15556_/X sky130_fd_sc_hd__buf_2
XANTENNA__16159__B1 _15761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12768_ _12765_/B _12767_/Y _12755_/X VGND VGND VPWR VPWR _12768_/X sky130_fd_sc_hd__and3_4
XPHY_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14507_ _14506_/X VGND VGND VPWR VPWR _14507_/Y sky130_fd_sc_hd__inv_2
X_11719_ _23802_/Q _11719_/B VGND VGND VPWR VPWR _11763_/A sky130_fd_sc_hd__or2_4
X_18275_ _18205_/A _18280_/B _18228_/X VGND VGND VPWR VPWR _18275_/Y sky130_fd_sc_hd__a21oi_4
X_15487_ _15472_/A VGND VGND VPWR VPWR _15487_/X sky130_fd_sc_hd__buf_2
X_12699_ _12638_/Y _12653_/X VGND VGND VPWR VPWR _12700_/B sky130_fd_sc_hd__or2_4
XANTENNA__18633__A _18633_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17226_ _11765_/X VGND VGND VPWR VPWR _17226_/X sky130_fd_sc_hd__buf_2
X_14438_ _24741_/Q VGND VGND VPWR VPWR _14541_/D sky130_fd_sc_hd__buf_2
XANTENNA__24455__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22155__A _22155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17157_ _17133_/A _17133_/B _17074_/A _17154_/Y VGND VGND VPWR VPWR _17157_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21455__B2 _21454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14369_ _14403_/A _14369_/B VGND VGND VPWR VPWR _14369_/X sky130_fd_sc_hd__or2_4
XANTENNA__16153__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16108_ _16107_/Y _16105_/X _15982_/X _16105_/X VGND VGND VPWR VPWR _24332_/D sky130_fd_sc_hd__a2bb2o_4
X_17088_ _17076_/X VGND VGND VPWR VPWR _17092_/B sky130_fd_sc_hd__inv_2
XANTENNA__16331__B1 _16254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16039_ _16038_/X VGND VGND VPWR VPWR _21882_/A sky130_fd_sc_hd__buf_2
XFILLER_130_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11728__C _11728_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22602__B _22524_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16634__B2 _16622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22707__A1 _22369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19729_ _21325_/B _19727_/X _19728_/X _19727_/X VGND VGND VPWR VPWR _19729_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18808__A _18807_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22740_ _23749_/Q _22173_/X _23717_/Q _22170_/X VGND VGND VPWR VPWR _22740_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_77_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22671_ _16336_/Y _21896_/X _16073_/Y _22549_/X VGND VGND VPWR VPWR _22671_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22049__B _13624_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21622_ _21625_/A _20043_/Y VGND VGND VPWR VPWR _21622_/X sky130_fd_sc_hd__or2_4
X_24410_ _24412_/CLK _15871_/X HRESETn VGND VGND VPWR VPWR _24410_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21553_ _21553_/A VGND VGND VPWR VPWR _21553_/X sky130_fd_sc_hd__buf_2
X_24341_ _23872_/CLK _16081_/X HRESETn VGND VGND VPWR VPWR _16080_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21888__B _22858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20504_ _22656_/A _20499_/X _20503_/Y VGND VGND VPWR VPWR _20504_/Y sky130_fd_sc_hd__a21oi_4
X_24272_ _24676_/CLK _16267_/X HRESETn VGND VGND VPWR VPWR _24272_/Q sky130_fd_sc_hd__dfrtp_4
X_21484_ _21169_/A _21484_/B VGND VGND VPWR VPWR _21484_/X sky130_fd_sc_hd__or2_4
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24196__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23223_ _23293_/CLK _23223_/D VGND VGND VPWR VPWR _23223_/Q sky130_fd_sc_hd__dfxtp_4
X_20435_ _15395_/Y _20416_/X _20425_/X _20434_/Y VGND VGND VPWR VPWR _20436_/A sky130_fd_sc_hd__o22a_4
XANTENNA__24125__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_210_0_HCLK clkbuf_8_211_0_HCLK/A VGND VGND VPWR VPWR _24201_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_107_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23154_ _23154_/CLK _23154_/D VGND VGND VPWR VPWR _23154_/Q sky130_fd_sc_hd__dfxtp_4
X_20366_ _20365_/X VGND VGND VPWR VPWR _23671_/D sky130_fd_sc_hd__inv_2
XANTENNA__16322__B1 _16153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22105_ _22105_/A _22101_/X _22104_/X VGND VGND VPWR VPWR _22105_/X sky130_fd_sc_hd__or3_4
X_23085_ _23085_/CLK _20118_/X VGND VGND VPWR VPWR _23085_/Q sky130_fd_sc_hd__dfxtp_4
X_20297_ _20297_/A _20293_/A VGND VGND VPWR VPWR _20297_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22512__B _22997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21749__A2 _21400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22946__A1 _21175_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22036_ _22036_/A VGND VGND VPWR VPWR _22246_/B sky130_fd_sc_hd__buf_2
XANTENNA__22946__B2 _22945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23781__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21128__B _21091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23760__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23987_ _23986_/CLK _23987_/D HRESETn VGND VGND VPWR VPWR _23987_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13740_ _13754_/A VGND VGND VPWR VPWR _13742_/B sky130_fd_sc_hd__inv_2
XFILLER_29_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17622__A _20778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22938_ _22997_/A _22938_/B _22931_/X _22937_/Y VGND VGND VPWR VPWR _22938_/X sky130_fd_sc_hd__or4_4
XFILLER_43_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21144__A _21144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13671_ _13647_/Y VGND VGND VPWR VPWR _13671_/X sky130_fd_sc_hd__buf_2
XFILLER_73_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24966__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22869_ _16490_/Y _22933_/B VGND VGND VPWR VPWR _22869_/X sky130_fd_sc_hd__and2_4
X_15410_ _22024_/B VGND VGND VPWR VPWR _15410_/X sky130_fd_sc_hd__buf_2
X_12622_ _12613_/X _12616_/X _12622_/C _12622_/D VGND VGND VPWR VPWR _12632_/C sky130_fd_sc_hd__or4_4
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24608_ _24182_/CLK _15343_/X HRESETn VGND VGND VPWR VPWR _24608_/Q sky130_fd_sc_hd__dfrtp_4
X_16390_ _11527_/Y VGND VGND VPWR VPWR _21109_/B sky130_fd_sc_hd__buf_2
XFILLER_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17060__C _17022_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20983__A _20961_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16074__A1_N _16073_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15341_ _22810_/A _15340_/X _11548_/X _15340_/X VGND VGND VPWR VPWR _24609_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ _25053_/Q VGND VGND VPWR VPWR _12553_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11622__B1 _11620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22882__B1 _20780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24539_ _23179_/CLK _24539_/D HRESETn VGND VGND VPWR VPWR _19821_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11504_ _21298_/B VGND VGND VPWR VPWR _16475_/A sky130_fd_sc_hd__buf_2
X_18060_ _18060_/A _18046_/X _18058_/X _18059_/X VGND VGND VPWR VPWR _18060_/X sky130_fd_sc_hd__or4_4
Xclkbuf_6_20_0_HCLK clkbuf_6_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_41_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15272_ _15285_/A VGND VGND VPWR VPWR _15272_/X sky130_fd_sc_hd__buf_2
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ _12474_/C _12466_/B _12453_/X _12481_/Y VGND VGND VPWR VPWR _12485_/A sky130_fd_sc_hd__a211o_4
XFILLER_138_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17011_ _16162_/A _17076_/A _16167_/Y _24047_/Q VGND VGND VPWR VPWR _17012_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13375__B1 _11631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14223_ _14223_/A VGND VGND VPWR VPWR _14223_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21437__A1 _24128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17069__A _24054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14154_ _18111_/B _14153_/X _14145_/X VGND VGND VPWR VPWR _24837_/D sky130_fd_sc_hd__a21o_4
X_13105_ _13016_/A VGND VGND VPWR VPWR _13309_/A sky130_fd_sc_hd__buf_2
XFILLER_98_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14085_ _14083_/Y _14079_/X _13668_/X _14084_/X VGND VGND VPWR VPWR _14085_/X sky130_fd_sc_hd__a2bb2o_4
X_18962_ _18961_/Y _18958_/X _18938_/X _18958_/X VGND VGND VPWR VPWR _23504_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23848__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13036_ _13011_/X _13027_/X _13035_/X VGND VGND VPWR VPWR _13036_/X sky130_fd_sc_hd__or3_4
X_17913_ _17817_/A _23144_/Q VGND VGND VPWR VPWR _17914_/C sky130_fd_sc_hd__or2_4
X_18893_ _18893_/A VGND VGND VPWR VPWR _18893_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15419__A2 _15415_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17844_ _17708_/X _17843_/X _23930_/Q _17767_/X VGND VGND VPWR VPWR _23930_/D sky130_fd_sc_hd__o22a_4
XFILLER_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17775_ _17881_/A _23148_/Q VGND VGND VPWR VPWR _17776_/C sky130_fd_sc_hd__or2_4
X_14987_ _14987_/A _15094_/A VGND VGND VPWR VPWR _14990_/B sky130_fd_sc_hd__or2_4
XANTENNA__12102__B2 _12101_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16726_ _16719_/X _16726_/B _16726_/C _16725_/X VGND VGND VPWR VPWR _16745_/A sky130_fd_sc_hd__or4_4
X_19514_ _19513_/Y _19511_/X _19445_/X _19511_/X VGND VGND VPWR VPWR _23309_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17532__A _17502_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13938_ _13936_/A VGND VGND VPWR VPWR _13938_/X sky130_fd_sc_hd__buf_2
XANTENNA__21373__B1 _21231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19445_ _19445_/A VGND VGND VPWR VPWR _19445_/X sky130_fd_sc_hd__buf_2
XANTENNA__21054__A _22249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16657_ _16652_/X _16653_/X _16096_/A _24105_/Q _16647_/X VGND VGND VPWR VPWR _24105_/D
+ sky130_fd_sc_hd__a32o_4
X_13869_ _13869_/A _13869_/B _24904_/Q _13869_/D VGND VGND VPWR VPWR _13870_/A sky130_fd_sc_hd__or4_4
Xclkbuf_7_102_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_205_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11580__A HWDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15608_ _12566_/Y _15604_/X _11566_/X _15607_/X VGND VGND VPWR VPWR _15608_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15052__A _24695_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19376_ _19375_/Y _19373_/X _19308_/X _19373_/X VGND VGND VPWR VPWR _23357_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16588_ _14860_/Y _16584_/X _16259_/X _16587_/X VGND VGND VPWR VPWR _16588_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21125__B1 _24396_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24636__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18327_ _18327_/A _18327_/B VGND VGND VPWR VPWR _18327_/X sky130_fd_sc_hd__or2_4
X_15539_ _19818_/A VGND VGND VPWR VPWR _19445_/A sky130_fd_sc_hd__buf_2
XFILLER_128_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19459__A _15556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11613__B1 _11612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18258_ _18258_/A _18459_/A VGND VGND VPWR VPWR _18258_/X sky130_fd_sc_hd__and2_4
XFILLER_72_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16552__B1 _16291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17209_ _17208_/Y _17206_/X _16546_/X _17206_/X VGND VGND VPWR VPWR _24016_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22625__B1 _22322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18189_ _21858_/A _23851_/Q _16119_/Y _18211_/A VGND VGND VPWR VPWR _18189_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20220_ _20232_/C VGND VGND VPWR VPWR _20220_/Y sky130_fd_sc_hd__inv_2
X_20151_ _20150_/Y _20148_/X _19963_/X _20148_/X VGND VGND VPWR VPWR _20151_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14935__A2_N _14933_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_40_0_HCLK clkbuf_7_20_0_HCLK/X VGND VGND VPWR VPWR _23514_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21229__A _21229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20082_ _20076_/Y VGND VGND VPWR VPWR _20082_/X sky130_fd_sc_hd__buf_2
XANTENNA__20133__A _23076_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23910_ _23908_/CLK _23910_/D HRESETn VGND VGND VPWR VPWR _23910_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14131__A _13492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24890_ _24783_/CLK _13972_/X HRESETn VGND VGND VPWR VPWR _24890_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23841_ _23824_/CLK _18458_/Y HRESETn VGND VGND VPWR VPWR _23841_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_61_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22156__A2 _15572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20984_ _20979_/A _20984_/B VGND VGND VPWR VPWR _20984_/X sky130_fd_sc_hd__or2_4
X_23772_ _24644_/CLK _20230_/X HRESETn VGND VGND VPWR VPWR _23772_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21364__B1 _20745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22723_ _12845_/Y _20838_/X _17502_/B _22191_/X VGND VGND VPWR VPWR _22723_/X sky130_fd_sc_hd__o22a_4
XFILLER_26_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19309__B1 _19308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24377__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22654_ _21850_/A VGND VGND VPWR VPWR _22654_/X sky130_fd_sc_hd__buf_2
XANTENNA__18178__A1_N _16068_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21605_ _21625_/A _21605_/B VGND VGND VPWR VPWR _21605_/X sky130_fd_sc_hd__or2_4
XANTENNA__15897__A _16376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24306__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22585_ _22585_/A VGND VGND VPWR VPWR _22585_/X sky130_fd_sc_hd__buf_2
XFILLER_22_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24324_ _24013_/CLK _24324_/D HRESETn VGND VGND VPWR VPWR _24324_/Q sky130_fd_sc_hd__dfrtp_4
X_21536_ _21535_/X VGND VGND VPWR VPWR _21536_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16543__B1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21411__B _21043_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21467_ _21333_/A _19677_/Y VGND VGND VPWR VPWR _21468_/C sky130_fd_sc_hd__or2_4
X_24255_ _24262_/CLK _24255_/D HRESETn VGND VGND VPWR VPWR _24255_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20418_ _20425_/A VGND VGND VPWR VPWR _20511_/A sky130_fd_sc_hd__buf_2
X_23206_ _23990_/CLK _19803_/X VGND VGND VPWR VPWR _23206_/Q sky130_fd_sc_hd__dfxtp_4
X_21398_ _23393_/Q _14016_/A _19225_/A _22042_/B VGND VGND VPWR VPWR _21398_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24186_ _24185_/CLK _16487_/X HRESETn VGND VGND VPWR VPWR _16485_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15649__A2 _15647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20349_ _17187_/A VGND VGND VPWR VPWR _20349_/X sky130_fd_sc_hd__buf_2
XFILLER_108_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23137_ _25106_/CLK _19983_/X VGND VGND VPWR VPWR _19981_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__23941__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25165__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21139__A _21333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23068_ _24112_/CLK HSEL VGND VGND VPWR VPWR _23032_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_95_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12155__A2_N _24575_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14910_ _24263_/Q VGND VGND VPWR VPWR _14910_/Y sky130_fd_sc_hd__inv_2
X_22019_ _21719_/A _22018_/X _16608_/Y _21408_/B VGND VGND VPWR VPWR _22019_/X sky130_fd_sc_hd__o22a_4
XFILLER_27_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15890_ _16369_/A VGND VGND VPWR VPWR _15890_/X sky130_fd_sc_hd__buf_2
X_14841_ _14832_/X _14834_/X _14837_/X _14840_/X VGND VGND VPWR VPWR _14841_/X sky130_fd_sc_hd__or4_4
XFILLER_76_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17560_ _16708_/Y _17564_/B _17559_/Y VGND VGND VPWR VPWR _17560_/X sky130_fd_sc_hd__o21a_4
X_14772_ _15045_/A _16649_/A _14770_/Y _16649_/A VGND VGND VPWR VPWR _14772_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11984_ _11983_/Y _11978_/X _11643_/X _11965_/Y VGND VGND VPWR VPWR _25148_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16511_ _16499_/A VGND VGND VPWR VPWR _16511_/X sky130_fd_sc_hd__buf_2
X_13723_ _13722_/X VGND VGND VPWR VPWR _13745_/A sky130_fd_sc_hd__inv_2
X_17491_ _16712_/Y _16700_/A _16685_/Y _17491_/D VGND VGND VPWR VPWR _17492_/D sky130_fd_sc_hd__or4_4
XFILLER_72_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19230_ _21252_/A _19226_/X _19207_/X _19226_/X VGND VGND VPWR VPWR _19230_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16442_ _16441_/Y _16439_/X _16093_/X _16439_/X VGND VGND VPWR VPWR _16442_/X sky130_fd_sc_hd__a2bb2o_4
X_13654_ _22355_/A _13652_/X _11594_/X _13652_/X VGND VGND VPWR VPWR _24937_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12605_ _12605_/A VGND VGND VPWR VPWR _12605_/Y sky130_fd_sc_hd__inv_2
X_19161_ _19159_/Y _19160_/X _19115_/X _19160_/X VGND VGND VPWR VPWR _23433_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16373_ _16373_/A VGND VGND VPWR VPWR _16373_/X sky130_fd_sc_hd__buf_2
XANTENNA__24047__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13585_ _13585_/A _13562_/B VGND VGND VPWR VPWR _13585_/Y sky130_fd_sc_hd__nand2_4
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18112_ _18112_/A VGND VGND VPWR VPWR _18118_/A sky130_fd_sc_hd__inv_2
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15324_ _24614_/Q VGND VGND VPWR VPWR _15324_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15600__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12536_ _12536_/A _12536_/B VGND VGND VPWR VPWR _12537_/C sky130_fd_sc_hd__nand2_4
X_19092_ _19078_/Y VGND VGND VPWR VPWR _19092_/X sky130_fd_sc_hd__buf_2
XFILLER_40_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12943__B _12947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18043_ _18043_/A VGND VGND VPWR VPWR _21147_/A sky130_fd_sc_hd__buf_2
XFILLER_129_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15255_ _13769_/B _15247_/X _15240_/X _13769_/A _15254_/X VGND VGND VPWR VPWR _24644_/D
+ sky130_fd_sc_hd__a32o_4
X_12467_ _12385_/Y _12467_/B VGND VGND VPWR VPWR _12468_/A sky130_fd_sc_hd__or2_4
XFILLER_8_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14206_ _14206_/A VGND VGND VPWR VPWR _20188_/A sky130_fd_sc_hd__inv_2
XFILLER_137_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15186_ _15158_/A VGND VGND VPWR VPWR _15192_/A sky130_fd_sc_hd__buf_2
XFILLER_126_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12398_ _12398_/A _12397_/X VGND VGND VPWR VPWR _12399_/A sky130_fd_sc_hd__or2_4
X_14137_ _24844_/Q _14120_/B _24843_/Q _14115_/X VGND VGND VPWR VPWR _14137_/X sky130_fd_sc_hd__o22a_4
X_19994_ _19993_/Y _19991_/X _19421_/X _19991_/X VGND VGND VPWR VPWR _19994_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23682__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_27_0_HCLK clkbuf_7_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_14068_ _13744_/X _14067_/X VGND VGND VPWR VPWR _14068_/X sky130_fd_sc_hd__or2_4
X_18945_ _18958_/A VGND VGND VPWR VPWR _18945_/X sky130_fd_sc_hd__buf_2
XFILLER_84_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12323__B2 _20808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13019_ _11732_/A VGND VGND VPWR VPWR _13075_/A sky130_fd_sc_hd__inv_2
X_18876_ _18875_/X VGND VGND VPWR VPWR _18876_/Y sky130_fd_sc_hd__inv_2
X_17827_ _17894_/A _17827_/B _17826_/X VGND VGND VPWR VPWR _17831_/B sky130_fd_sc_hd__and3_4
XANTENNA__24888__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15273__B1 _14228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17758_ _17961_/A _17755_/X _17757_/X VGND VGND VPWR VPWR _17758_/X sky130_fd_sc_hd__and3_4
XANTENNA__24817__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17014__B2 _17021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16709_ _22639_/A _23961_/Q _15952_/Y _16708_/Y VGND VGND VPWR VPWR _16709_/X sky130_fd_sc_hd__o22a_4
X_17689_ _16022_/Y VGND VGND VPWR VPWR _17689_/X sky130_fd_sc_hd__buf_2
XFILLER_120_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19428_ _19427_/Y _19425_/X _19381_/X _19425_/X VGND VGND VPWR VPWR _23339_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24470__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22608__A _13334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19359_ _13210_/B VGND VGND VPWR VPWR _19359_/Y sky130_fd_sc_hd__inv_2
X_22370_ _16188_/A _21984_/X VGND VGND VPWR VPWR _22370_/X sky130_fd_sc_hd__or2_4
X_21321_ _21079_/X _21318_/Y _13334_/X _21320_/X VGND VGND VPWR VPWR _21322_/A sky130_fd_sc_hd__o22a_4
XFILLER_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21252_ _21252_/A _20827_/X VGND VGND VPWR VPWR _21252_/X sky130_fd_sc_hd__or2_4
X_24040_ _24606_/CLK _17129_/X HRESETn VGND VGND VPWR VPWR _24040_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14551__A2 _14437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20203_ _23771_/Q VGND VGND VPWR VPWR _20203_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21183_ _11941_/X _21181_/X _21182_/X _18013_/Y _21716_/B VGND VGND VPWR VPWR _21184_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_137_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20134_ _11734_/Y _11746_/Y _20134_/C VGND VGND VPWR VPWR _20134_/X sky130_fd_sc_hd__or3_4
X_20065_ _20054_/X _15410_/X _18000_/X _20064_/X _20055_/X VGND VGND VPWR VPWR _23105_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_86_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14889__A2_N _14887_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19652__A _19646_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24942_ _24944_/CLK _13642_/X HRESETn VGND VGND VPWR VPWR _24942_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20798__A _22870_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24873_ _23657_/CLK _14042_/X HRESETn VGND VGND VPWR VPWR _14041_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23824_ _23824_/CLK _23824_/D HRESETn VGND VGND VPWR VPWR _18420_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24558__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23755_ _24185_/CLK _23755_/D HRESETn VGND VGND VPWR VPWR _23755_/Q sky130_fd_sc_hd__dfrtp_4
X_20967_ _20967_/A _20967_/B _20967_/C VGND VGND VPWR VPWR _20967_/X sky130_fd_sc_hd__and3_4
X_22706_ _22706_/A _22638_/X VGND VGND VPWR VPWR _22706_/X sky130_fd_sc_hd__or2_4
X_23686_ _23664_/CLK _23686_/D HRESETn VGND VGND VPWR VPWR _14633_/A sky130_fd_sc_hd__dfrtp_4
X_20898_ _20836_/X _20840_/X _20897_/Y VGND VGND VPWR VPWR _20898_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21422__A _16041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24140__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22637_ _22637_/A VGND VGND VPWR VPWR _22637_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15420__A _22314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13370_ _13370_/A VGND VGND VPWR VPWR _13370_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16516__B1 _16179_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20312__A1 _14259_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22568_ _16513_/Y _22011_/A _15361_/Y _22452_/X VGND VGND VPWR VPWR _22568_/X sky130_fd_sc_hd__o22a_4
XFILLER_10_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16235__B _16235_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12321_ _12469_/A _12319_/Y _25097_/Q _12320_/Y VGND VGND VPWR VPWR _12321_/X sky130_fd_sc_hd__a2bb2o_4
X_24307_ _24307_/CLK _24307_/D HRESETn VGND VGND VPWR VPWR _16172_/A sky130_fd_sc_hd__dfrtp_4
X_21519_ _21519_/A _21519_/B _21518_/X VGND VGND VPWR VPWR _21519_/X sky130_fd_sc_hd__and3_4
XFILLER_10_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22499_ _21870_/A _22497_/X _21886_/X _22498_/X VGND VGND VPWR VPWR _22499_/X sky130_fd_sc_hd__o22a_4
X_15040_ _15033_/A _15020_/X _15027_/X _15038_/B VGND VGND VPWR VPWR _15041_/A sky130_fd_sc_hd__a211o_4
X_12252_ _12227_/X _12252_/B _12251_/X VGND VGND VPWR VPWR _25117_/D sky130_fd_sc_hd__and3_4
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24238_ _24244_/CLK _16348_/X HRESETn VGND VGND VPWR VPWR _16345_/A sky130_fd_sc_hd__dfrtp_4
X_12183_ _12183_/A _12183_/B VGND VGND VPWR VPWR _12184_/D sky130_fd_sc_hd__or2_4
XFILLER_134_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24169_ _24168_/CLK _16528_/X HRESETn VGND VGND VPWR VPWR _16527_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16251__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23014__B1 _24058_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16991_ _16964_/X _16972_/X _16981_/X _16991_/D VGND VGND VPWR VPWR _16991_/X sky130_fd_sc_hd__or4_4
XFILLER_27_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15942_ _15940_/Y _15936_/X _15761_/X _15941_/X VGND VGND VPWR VPWR _15942_/X sky130_fd_sc_hd__a2bb2o_4
X_18730_ _17952_/B VGND VGND VPWR VPWR _18730_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18661_ _18661_/A VGND VGND VPWR VPWR _21001_/B sky130_fd_sc_hd__inv_2
X_15873_ _15885_/A VGND VGND VPWR VPWR _15873_/X sky130_fd_sc_hd__buf_2
XFILLER_37_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24981__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16598__A3 _11585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14824_ _14997_/A _14823_/Y _15092_/A _24126_/Q VGND VGND VPWR VPWR _14829_/B sky130_fd_sc_hd__a2bb2o_4
X_17612_ _17611_/X VGND VGND VPWR VPWR _23946_/D sky130_fd_sc_hd__inv_2
XFILLER_76_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17082__A _17052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18592_ _18592_/A _18592_/B _18590_/X _18591_/X VGND VGND VPWR VPWR _18592_/X sky130_fd_sc_hd__or4_4
XANTENNA__24299__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24910__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17543_ _17509_/A _17534_/B _17542_/X VGND VGND VPWR VPWR _23965_/D sky130_fd_sc_hd__and3_4
X_14755_ _24098_/Q VGND VGND VPWR VPWR _14755_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24228__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11967_ _11959_/Y _11966_/X _11612_/X _11966_/X VGND VGND VPWR VPWR _25155_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22540__A2 _22539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18906__A _18899_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13706_ _24915_/Q _13686_/X _24914_/Q _13681_/X VGND VGND VPWR VPWR _13706_/X sky130_fd_sc_hd__o22a_4
X_17474_ _21801_/A VGND VGND VPWR VPWR _17474_/Y sky130_fd_sc_hd__inv_2
X_14686_ _14686_/A VGND VGND VPWR VPWR _24717_/D sky130_fd_sc_hd__inv_2
X_11898_ _11884_/B VGND VGND VPWR VPWR _11898_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22428__A _21434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16425_ _24209_/Q VGND VGND VPWR VPWR _16425_/Y sky130_fd_sc_hd__inv_2
X_19213_ _19212_/Y VGND VGND VPWR VPWR _19213_/X sky130_fd_sc_hd__buf_2
XANTENNA__21332__A _21469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13637_ _13637_/A VGND VGND VPWR VPWR _13637_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16426__A _16426_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19144_ _19144_/A _19144_/B _18874_/X VGND VGND VPWR VPWR _19144_/X sky130_fd_sc_hd__or3_4
X_16356_ _24234_/Q VGND VGND VPWR VPWR _16356_/Y sky130_fd_sc_hd__inv_2
X_13568_ _23904_/Q _13568_/B VGND VGND VPWR VPWR _13568_/X sky130_fd_sc_hd__and2_4
XANTENNA__16507__B1 _16259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15307_ _16038_/B _15304_/X HADDR[20] _15304_/X VGND VGND VPWR VPWR _15307_/X sky130_fd_sc_hd__a2bb2o_4
X_12519_ _12509_/A _12515_/X _12519_/C VGND VGND VPWR VPWR _12519_/X sky130_fd_sc_hd__and3_4
X_19075_ _19075_/A VGND VGND VPWR VPWR _19075_/Y sky130_fd_sc_hd__inv_2
X_16287_ _14937_/Y _16286_/X _15897_/X _16286_/X VGND VGND VPWR VPWR _16287_/X sky130_fd_sc_hd__a2bb2o_4
X_13499_ _13499_/A _21020_/A VGND VGND VPWR VPWR _13499_/Y sky130_fd_sc_hd__nor2_4
XFILLER_117_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23863__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18026_ _23903_/Q VGND VGND VPWR VPWR _19530_/A sky130_fd_sc_hd__inv_2
X_15238_ _23685_/Q _14072_/A _14071_/D _15237_/X VGND VGND VPWR VPWR _15241_/A sky130_fd_sc_hd__o22a_4
XANTENNA__25087__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22163__A _22163_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25016__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15169_ _14950_/Y _15168_/X VGND VGND VPWR VPWR _15183_/B sky130_fd_sc_hd__or2_4
XFILLER_114_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18680__B1 _18679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19977_ _19977_/A VGND VGND VPWR VPWR _19977_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18928_ _18926_/Y _18922_/X _18883_/X _18927_/X VGND VGND VPWR VPWR _23516_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18859_ _18854_/A VGND VGND VPWR VPWR _18859_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_114_0_HCLK clkbuf_7_57_0_HCLK/X VGND VGND VPWR VPWR _24923_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16589__A3 HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15505__A HWDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_177_0_HCLK clkbuf_7_88_0_HCLK/X VGND VGND VPWR VPWR _25021_/CLK sky130_fd_sc_hd__clkbuf_1
X_21870_ _21870_/A _21870_/B VGND VGND VPWR VPWR _21870_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__21319__B1 _12818_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24651__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20790__B2 _15637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20821_ _22148_/A VGND VGND VPWR VPWR _20821_/X sky130_fd_sc_hd__buf_2
XFILLER_78_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23540_ _23133_/CLK _18860_/X VGND VGND VPWR VPWR _23540_/Q sky130_fd_sc_hd__dfxtp_4
X_20752_ _20751_/X VGND VGND VPWR VPWR _20753_/A sky130_fd_sc_hd__buf_2
XFILLER_126_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23685__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24771__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20683_ _20550_/A _23758_/Q _13543_/B _24189_/Q _20602_/X VGND VGND VPWR VPWR _20683_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_91_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23471_ _23471_/CLK _19054_/X VGND VGND VPWR VPWR _13308_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25210_ _25214_/CLK _11564_/X HRESETn VGND VGND VPWR VPWR _11562_/A sky130_fd_sc_hd__dfrtp_4
X_22422_ _22418_/X _22419_/X _22421_/X VGND VGND VPWR VPWR _22457_/A sky130_fd_sc_hd__and3_4
XANTENNA__21098__A2 _21097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25141_ _25141_/CLK _25141_/D HRESETn VGND VGND VPWR VPWR _12004_/A sky130_fd_sc_hd__dfrtp_4
X_22353_ _24234_/Q _22147_/X _20799_/X _22352_/X VGND VGND VPWR VPWR _22353_/X sky130_fd_sc_hd__a211o_4
XANTENNA__19647__A _19646_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21304_ _12006_/Y _13357_/X _18124_/Y _21083_/X VGND VGND VPWR VPWR _21304_/X sky130_fd_sc_hd__o22a_4
X_22284_ _22500_/A _22284_/B VGND VGND VPWR VPWR _22292_/C sky130_fd_sc_hd__nor2_4
X_25072_ _25091_/CLK _25072_/D HRESETn VGND VGND VPWR VPWR _12348_/A sky130_fd_sc_hd__dfrtp_4
X_21235_ _21235_/A _21235_/B VGND VGND VPWR VPWR _21235_/X sky130_fd_sc_hd__or2_4
XANTENNA__19999__B1 _15520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24023_ _23664_/CLK _24023_/D HRESETn VGND VGND VPWR VPWR _20723_/A sky130_fd_sc_hd__dfstp_4
XFILLER_105_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17167__A _17086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16277__A2 _16276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21166_ _21935_/A _21166_/B VGND VGND VPWR VPWR _21166_/X sky130_fd_sc_hd__or2_4
XFILLER_46_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18671__B1 _17202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22801__A _22777_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15485__B1 _24568_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20117_ _20116_/X VGND VGND VPWR VPWR _20117_/X sky130_fd_sc_hd__buf_2
XFILLER_120_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_10_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21097_ _21097_/A _21097_/B VGND VGND VPWR VPWR _21097_/X sky130_fd_sc_hd__and2_4
XFILLER_59_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12104__A _24552_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24739__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_73_0_HCLK clkbuf_7_73_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_73_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20048_ _20035_/Y VGND VGND VPWR VPWR _20048_/X sky130_fd_sc_hd__buf_2
X_24925_ _24937_/CLK _24925_/D HRESETn VGND VGND VPWR VPWR _24925_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21310__A2_N _20826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11943__A _22616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15415__A _16475_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12870_ _12812_/Y _12899_/C VGND VGND VPWR VPWR _12894_/A sky130_fd_sc_hd__or2_4
XFILLER_46_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24392__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24856_ _23657_/CLK _14095_/X HRESETn VGND VGND VPWR VPWR _24856_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11821_ _11817_/A _11823_/A VGND VGND VPWR VPWR _11821_/Y sky130_fd_sc_hd__nor2_4
X_23807_ _23648_/CLK _18629_/X HRESETn VGND VGND VPWR VPWR _23807_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_61_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24321__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24787_ _24788_/CLK _14298_/X HRESETn VGND VGND VPWR VPWR _14297_/A sky130_fd_sc_hd__dfrtp_4
X_21999_ _16685_/A _21850_/A VGND VGND VPWR VPWR _21999_/X sky130_fd_sc_hd__and2_4
XFILLER_14_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14539_/Y VGND VGND VPWR VPWR _14540_/X sky130_fd_sc_hd__buf_2
XPHY_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11751_/X VGND VGND VPWR VPWR _11753_/A sky130_fd_sc_hd__buf_2
XFILLER_121_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23738_ _24259_/CLK _20608_/X HRESETn VGND VGND VPWR VPWR _23738_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14471_/A VGND VGND VPWR VPWR _14471_/X sky130_fd_sc_hd__buf_2
XFILLER_70_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11683_/A VGND VGND VPWR VPWR _11683_/Y sky130_fd_sc_hd__inv_2
XPHY_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23669_ _24723_/CLK _23669_/D HRESETn VGND VGND VPWR VPWR _17173_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16246__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _24292_/Q VGND VGND VPWR VPWR _16210_/Y sky130_fd_sc_hd__inv_2
XPHY_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _13421_/Y _14424_/A _13421_/Y _14424_/A VGND VGND VPWR VPWR _13422_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17190_ _17171_/X _17185_/X _24024_/Q _24025_/Q _17188_/X VGND VGND VPWR VPWR _24025_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22286__B2 _22285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16141_ HWDATA[30] VGND VGND VPWR VPWR _16141_/X sky130_fd_sc_hd__buf_2
X_13353_ _13353_/A VGND VGND VPWR VPWR _13353_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17162__B1 _17057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12304_ _12508_/A _24478_/Q _12508_/A _24478_/Q VGND VGND VPWR VPWR _12312_/A sky130_fd_sc_hd__a2bb2o_4
X_16072_ _16070_/Y _16071_/X _15855_/X _16071_/X VGND VGND VPWR VPWR _16072_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22038__B2 _20866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25180__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13284_ _13316_/A _13284_/B VGND VGND VPWR VPWR _13284_/X sky130_fd_sc_hd__or2_4
X_15023_ _15025_/B VGND VGND VPWR VPWR _15023_/Y sky130_fd_sc_hd__inv_2
X_19900_ _21221_/B _19897_/X _19835_/X _19897_/X VGND VGND VPWR VPWR _19900_/X sky130_fd_sc_hd__a2bb2o_4
X_12235_ _12149_/Y _12229_/X _12203_/X _12232_/B VGND VGND VPWR VPWR _12235_/X sky130_fd_sc_hd__a211o_4
XANTENNA__14704__A2_N _24118_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19831_ _19831_/A VGND VGND VPWR VPWR _19831_/X sky130_fd_sc_hd__buf_2
X_12166_ _12165_/X VGND VGND VPWR VPWR _12190_/A sky130_fd_sc_hd__buf_2
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15476__B1 _11540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19762_ _23221_/Q VGND VGND VPWR VPWR _19762_/Y sky130_fd_sc_hd__inv_2
X_12097_ _12097_/A VGND VGND VPWR VPWR _12097_/Y sky130_fd_sc_hd__inv_2
X_16974_ _16172_/A _24045_/Q _16172_/Y _17042_/A VGND VGND VPWR VPWR _16981_/A sky130_fd_sc_hd__o22a_4
X_18713_ _18710_/Y _18705_/X _18712_/X _18697_/A VGND VGND VPWR VPWR _18713_/X sky130_fd_sc_hd__a2bb2o_4
X_15925_ _24390_/Q VGND VGND VPWR VPWR _15925_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19693_ _19693_/A VGND VGND VPWR VPWR _19693_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24409__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11853__A _19610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15856_ _15853_/Y _15854_/X _15855_/X _15854_/X VGND VGND VPWR VPWR _15856_/X sky130_fd_sc_hd__a2bb2o_4
X_18644_ _18644_/A VGND VGND VPWR VPWR _18644_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14261__A1_N _14259_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14807_ _15085_/A _24125_/Q _15085_/A _24125_/Q VGND VGND VPWR VPWR _14807_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24062__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15787_ _15767_/X VGND VGND VPWR VPWR _15787_/X sky130_fd_sc_hd__buf_2
X_18575_ _16383_/A _23815_/Q _16383_/Y _18552_/A VGND VGND VPWR VPWR _18575_/X sky130_fd_sc_hd__o22a_4
X_12999_ _12999_/A _13008_/B VGND VGND VPWR VPWR _12999_/X sky130_fd_sc_hd__or2_4
XFILLER_79_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18636__A _21188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19914__B1 _19825_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14738_ _24701_/Q _14737_/A _14736_/X _14737_/Y VGND VGND VPWR VPWR _14749_/A sky130_fd_sc_hd__o22a_4
X_17526_ _17515_/D _17524_/A VGND VGND VPWR VPWR _17526_/X sky130_fd_sc_hd__or2_4
XFILLER_75_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21721__B1 _14801_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22158__A _21050_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21062__A _20820_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17457_ _21801_/A _17457_/B VGND VGND VPWR VPWR _17457_/Y sky130_fd_sc_hd__nand2_4
X_14669_ _14655_/X _14668_/Y _24721_/Q _14655_/X VGND VGND VPWR VPWR _14669_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16408_ _24216_/Q VGND VGND VPWR VPWR _16408_/Y sky130_fd_sc_hd__inv_2
X_17388_ _17390_/A _17382_/X _17388_/C VGND VGND VPWR VPWR _17388_/X sky130_fd_sc_hd__and3_4
X_16339_ _16339_/A VGND VGND VPWR VPWR _16339_/X sky130_fd_sc_hd__buf_2
X_19127_ _17714_/B VGND VGND VPWR VPWR _19127_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19058_ _19071_/A VGND VGND VPWR VPWR _19058_/X sky130_fd_sc_hd__buf_2
XFILLER_106_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12517__A1 _12345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18009_ _18005_/Y _18008_/X _16546_/X _18008_/X VGND VGND VPWR VPWR _23909_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21020_ _21020_/A _21020_/B VGND VGND VPWR VPWR _21020_/X sky130_fd_sc_hd__and2_4
XFILLER_86_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15467__B1 _24576_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24832__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22971_ _22971_/A _22970_/X VGND VGND VPWR VPWR _22971_/X sky130_fd_sc_hd__and2_4
XFILLER_68_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14229__A1_N _14223_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24710_ _24674_/CLK _24710_/D HRESETn VGND VGND VPWR VPWR _24710_/Q sky130_fd_sc_hd__dfrtp_4
X_21922_ _20968_/X _21918_/X _21921_/X VGND VGND VPWR VPWR _21922_/X sky130_fd_sc_hd__or3_4
XFILLER_55_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24641_ _24641_/CLK _15259_/X HRESETn VGND VGND VPWR VPWR _13716_/D sky130_fd_sc_hd__dfrtp_4
X_21853_ _20783_/X _21851_/X _22629_/A _12596_/A _21047_/A VGND VGND VPWR VPWR _21853_/X
+ sky130_fd_sc_hd__a32o_4
X_20804_ _22014_/B _20803_/X _24499_/Q _21591_/B VGND VGND VPWR VPWR _20804_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20674__A1_N _20556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24572_ _24573_/CLK _24572_/D HRESETn VGND VGND VPWR VPWR _12089_/A sky130_fd_sc_hd__dfrtp_4
X_21784_ _21760_/X _21784_/B VGND VGND VPWR VPWR _21784_/X sky130_fd_sc_hd__or2_4
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23523_ _23531_/CLK _23523_/D VGND VGND VPWR VPWR _17834_/B sky130_fd_sc_hd__dfxtp_4
X_20735_ _20735_/A _20735_/B VGND VGND VPWR VPWR _20735_/X sky130_fd_sc_hd__and2_4
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16066__A _24347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23785__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22268__B2 _13619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22218__D _22510_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14745__A2 _14744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23454_ _24735_/CLK _19102_/X VGND VGND VPWR VPWR _23454_/Q sky130_fd_sc_hd__dfxtp_4
X_20666_ _20647_/X _20665_/X _16492_/A _20651_/X VGND VGND VPWR VPWR _23752_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23714__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22405_ _11691_/Y _20902_/X _13450_/Y _20918_/X VGND VGND VPWR VPWR _22405_/X sky130_fd_sc_hd__o22a_4
X_20597_ _20597_/A VGND VGND VPWR VPWR _20597_/Y sky130_fd_sc_hd__inv_2
X_23385_ _23385_/CLK _19297_/X VGND VGND VPWR VPWR _19295_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24629__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25124_ _25130_/CLK _25124_/D HRESETn VGND VGND VPWR VPWR _25124_/Q sky130_fd_sc_hd__dfrtp_4
X_22336_ _24105_/Q _22574_/B VGND VGND VPWR VPWR _22341_/B sky130_fd_sc_hd__or2_4
XFILLER_125_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25055_ _24521_/CLK _25055_/D HRESETn VGND VGND VPWR VPWR _25055_/Q sky130_fd_sc_hd__dfrtp_4
X_22267_ _22267_/A _22314_/B VGND VGND VPWR VPWR _22267_/X sky130_fd_sc_hd__and2_4
XFILLER_133_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12020_ _12014_/B VGND VGND VPWR VPWR _12020_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24006_ _24005_/CLK _24006_/D HRESETn VGND VGND VPWR VPWR _24006_/Q sky130_fd_sc_hd__dfrtp_4
X_21218_ _14471_/X _21208_/X _21217_/X VGND VGND VPWR VPWR _21218_/X sky130_fd_sc_hd__or3_4
X_22198_ _22198_/A VGND VGND VPWR VPWR _22198_/X sky130_fd_sc_hd__buf_2
XFILLER_2_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22531__A _21069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20451__B1 _20446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22991__A2 _20926_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21149_ _21339_/A _21141_/X _21148_/X VGND VGND VPWR VPWR _21149_/X sky130_fd_sc_hd__or3_4
XANTENNA__24573__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22250__B _22999_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13971_ _13952_/A VGND VGND VPWR VPWR _13971_/X sky130_fd_sc_hd__buf_2
XFILLER_19_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24502__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15710_ _12356_/Y _15702_/X _15709_/X _15666_/A VGND VGND VPWR VPWR _24468_/D sky130_fd_sc_hd__a2bb2o_4
X_12922_ _12922_/A VGND VGND VPWR VPWR _12922_/X sky130_fd_sc_hd__buf_2
XFILLER_20_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24908_ _24904_/CLK _24908_/D HRESETn VGND VGND VPWR VPWR _13816_/A sky130_fd_sc_hd__dfrtp_4
X_16690_ _22256_/A VGND VGND VPWR VPWR _17490_/A sky130_fd_sc_hd__inv_2
X_15641_ _22218_/C VGND VGND VPWR VPWR _15641_/X sky130_fd_sc_hd__buf_2
XFILLER_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12853_ _12853_/A VGND VGND VPWR VPWR _12853_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_160_0_HCLK clkbuf_7_80_0_HCLK/X VGND VGND VPWR VPWR _23179_/CLK sky130_fd_sc_hd__clkbuf_1
X_24839_ _24840_/CLK _14148_/X HRESETn VGND VGND VPWR VPWR _24839_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_3_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11804_ _11804_/A VGND VGND VPWR VPWR _11804_/Y sky130_fd_sc_hd__inv_2
X_18360_ _23821_/Q VGND VGND VPWR VPWR _18361_/A sky130_fd_sc_hd__inv_2
X_15572_ _15572_/A VGND VGND VPWR VPWR _22223_/A sky130_fd_sc_hd__buf_2
XANTENNA__21894__A2_N _21544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_17_0_HCLK clkbuf_7_8_0_HCLK/X VGND VGND VPWR VPWR _24841_/CLK sky130_fd_sc_hd__clkbuf_1
X_12784_ _22527_/A VGND VGND VPWR VPWR _12785_/A sky130_fd_sc_hd__inv_2
XPHY_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17311_/A VGND VGND VPWR VPWR _17311_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14523_/A VGND VGND VPWR VPWR _14524_/D sky130_fd_sc_hd__buf_2
XPHY_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11735_ _23893_/Q VGND VGND VPWR VPWR _11735_/Y sky130_fd_sc_hd__inv_2
X_18291_ _18263_/A _18218_/C VGND VGND VPWR VPWR _18292_/B sky130_fd_sc_hd__or2_4
XPHY_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17383__B1 _17336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17236_/X _17238_/X _17242_/C _17241_/X VGND VGND VPWR VPWR _17269_/A sky130_fd_sc_hd__or4_4
XPHY_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _14528_/A VGND VGND VPWR VPWR _21010_/A sky130_fd_sc_hd__buf_2
XPHY_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _13549_/A _22484_/A _24958_/Q _22319_/A VGND VGND VPWR VPWR _11666_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _15712_/A _15713_/A VGND VGND VPWR VPWR _13471_/A sky130_fd_sc_hd__or2_4
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17173_ _17173_/A _17173_/B VGND VGND VPWR VPWR _17174_/B sky130_fd_sc_hd__or2_4
XANTENNA__20809__A2 _20805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14385_ _14385_/A _14384_/X VGND VGND VPWR VPWR _14386_/A sky130_fd_sc_hd__or2_4
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11597_ HWDATA[11] VGND VGND VPWR VPWR _16100_/A sky130_fd_sc_hd__buf_2
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16124_ _21097_/A _16046_/A _15709_/X _16046_/A VGND VGND VPWR VPWR _24325_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22425__B _22147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13336_ _13335_/X VGND VGND VPWR VPWR _13337_/A sky130_fd_sc_hd__buf_2
XANTENNA__15697__B1 _15511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16055_ _16054_/Y _16052_/X _15837_/X _16052_/X VGND VGND VPWR VPWR _24352_/D sky130_fd_sc_hd__a2bb2o_4
X_13267_ _13299_/A _13267_/B _13267_/C VGND VGND VPWR VPWR _13271_/B sky130_fd_sc_hd__and3_4
X_15006_ _15006_/A VGND VGND VPWR VPWR _15006_/Y sky130_fd_sc_hd__inv_2
X_12218_ _12079_/X _12216_/X _12217_/Y VGND VGND VPWR VPWR _25127_/D sky130_fd_sc_hd__o21a_4
XFILLER_29_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13198_ _13230_/A _20000_/A VGND VGND VPWR VPWR _13198_/X sky130_fd_sc_hd__or2_4
XANTENNA__22441__A _21572_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19814_ _19831_/A VGND VGND VPWR VPWR _19814_/X sky130_fd_sc_hd__buf_2
X_12149_ _25122_/Q VGND VGND VPWR VPWR _12149_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22160__B _22952_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21057__A _21432_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19745_ _23227_/Q VGND VGND VPWR VPWR _21629_/B sky130_fd_sc_hd__inv_2
X_16957_ _16837_/D _16879_/X _16858_/X _16954_/Y VGND VGND VPWR VPWR _16958_/A sky130_fd_sc_hd__a211o_4
XFILLER_81_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24243__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15908_ _24395_/Q VGND VGND VPWR VPWR _15908_/Y sky130_fd_sc_hd__inv_2
X_19676_ _19675_/Y _19673_/X _19607_/X _19673_/X VGND VGND VPWR VPWR _23251_/D sky130_fd_sc_hd__a2bb2o_4
X_16888_ _16760_/A _16888_/B VGND VGND VPWR VPWR _16888_/X sky130_fd_sc_hd__or2_4
XFILLER_53_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18627_ _18607_/X _18621_/X _23646_/Q _23809_/Q _18624_/X VGND VGND VPWR VPWR _18627_/X
+ sky130_fd_sc_hd__a32o_4
X_15839_ _24422_/Q VGND VGND VPWR VPWR _15839_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18558_ _18484_/A _18552_/B _18558_/C VGND VGND VPWR VPWR _18558_/X sky130_fd_sc_hd__and3_4
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18085__B _18080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17509_ _17509_/A _17509_/B _17509_/C VGND VGND VPWR VPWR _17509_/X sky130_fd_sc_hd__and3_4
X_18489_ _18491_/B VGND VGND VPWR VPWR _18489_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13303__A _13271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20520_ _20520_/A VGND VGND VPWR VPWR _20520_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14727__A2 _14726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22616__A _22616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20451_ _22008_/A _20437_/X _20446_/X _20450_/X VGND VGND VPWR VPWR _20451_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25031__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20382_ _20385_/B _20381_/Y _20373_/X VGND VGND VPWR VPWR _20382_/X sky130_fd_sc_hd__and3_4
X_23170_ _23308_/CLK _19895_/X VGND VGND VPWR VPWR _19894_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_101_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22121_ _21064_/Y VGND VGND VPWR VPWR _22121_/X sky130_fd_sc_hd__buf_2
XANTENNA__20681__B1 _13543_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22052_ _21667_/X _19009_/Y VGND VGND VPWR VPWR _22052_/X sky130_fd_sc_hd__or2_4
XFILLER_133_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22351__A _22351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21003_ _21010_/A _21001_/X _21003_/C VGND VGND VPWR VPWR _21003_/X sky130_fd_sc_hd__and3_4
XFILLER_87_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22954_ _24424_/Q _22281_/X _20782_/A _22953_/X VGND VGND VPWR VPWR _22955_/C sky130_fd_sc_hd__a211o_4
X_21905_ _21905_/A _21905_/B _21905_/C _21905_/D VGND VGND VPWR VPWR _21905_/X sky130_fd_sc_hd__or4_4
X_22885_ _21561_/X _22883_/X _21562_/X _22884_/X VGND VGND VPWR VPWR _22885_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23966__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_233_0_HCLK clkbuf_8_233_0_HCLK/A VGND VGND VPWR VPWR _24604_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22489__A1 _22322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24624_ _24643_/CLK _15293_/X HRESETn VGND VGND VPWR VPWR _24624_/Q sky130_fd_sc_hd__dfrtp_4
X_21836_ _17636_/A _21814_/Y _21821_/Y _21829_/Y _21835_/Y VGND VGND VPWR VPWR _21836_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_43_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25119__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24555_ _24566_/CLK _24555_/D HRESETn VGND VGND VPWR VPWR _24555_/Q sky130_fd_sc_hd__dfrtp_4
X_21767_ _21519_/A _21767_/B _21766_/X VGND VGND VPWR VPWR _21767_/X sky130_fd_sc_hd__and3_4
XFILLER_70_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ _11599_/A VGND VGND VPWR VPWR _11521_/A sky130_fd_sc_hd__buf_2
XANTENNA__13213__A _13309_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23506_ _23514_/CLK _18956_/X VGND VGND VPWR VPWR _17871_/B sky130_fd_sc_hd__dfxtp_4
X_20718_ _14012_/Y _23654_/Q _13800_/A VGND VGND VPWR VPWR _23654_/D sky130_fd_sc_hd__a21o_4
XFILLER_71_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24486_ _24488_/CLK _24486_/D HRESETn VGND VGND VPWR VPWR _24486_/Q sky130_fd_sc_hd__dfrtp_4
X_21698_ _21695_/X _21696_/X _21697_/X VGND VGND VPWR VPWR _21698_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23437_ _25067_/CLK _19150_/X VGND VGND VPWR VPWR _23437_/Q sky130_fd_sc_hd__dfxtp_4
X_20649_ _23748_/Q _13524_/B _20653_/A _13524_/D VGND VGND VPWR VPWR _20649_/X sky130_fd_sc_hd__or4_4
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14170_ _12053_/A _14170_/B _14170_/C VGND VGND VPWR VPWR _24833_/D sky130_fd_sc_hd__and3_4
X_23368_ _24998_/CLK _19344_/X VGND VGND VPWR VPWR _13273_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15679__B1 _11563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13121_ _13120_/X _23540_/Q VGND VGND VPWR VPWR _13121_/X sky130_fd_sc_hd__or2_4
X_25107_ _25123_/CLK _25107_/D HRESETn VGND VGND VPWR VPWR _12122_/A sky130_fd_sc_hd__dfrtp_4
X_22319_ _22319_/A _21180_/X VGND VGND VPWR VPWR _22319_/X sky130_fd_sc_hd__and2_4
XANTENNA__24754__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23299_ _23939_/CLK _19542_/X VGND VGND VPWR VPWR _23299_/Q sky130_fd_sc_hd__dfxtp_4
X_13052_ _13113_/A _13044_/X _13051_/X _11708_/A _11708_/B VGND VGND VPWR VPWR _13052_/X
+ sky130_fd_sc_hd__o32a_4
X_25038_ _25044_/CLK _25038_/D HRESETn VGND VGND VPWR VPWR _12650_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15694__A3 _16100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12003_ _12001_/Y _12002_/X _11626_/X _12002_/X VGND VGND VPWR VPWR _25142_/D sky130_fd_sc_hd__a2bb2o_4
X_17860_ _17924_/A _17860_/B VGND VGND VPWR VPWR _17862_/B sky130_fd_sc_hd__or2_4
XFILLER_120_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16811_ _16811_/A _16811_/B VGND VGND VPWR VPWR _17132_/A sky130_fd_sc_hd__or2_4
X_17791_ _17895_/A _23460_/Q VGND VGND VPWR VPWR _17791_/X sky130_fd_sc_hd__or2_4
XFILLER_94_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19530_ _19530_/A VGND VGND VPWR VPWR _19530_/X sky130_fd_sc_hd__buf_2
X_13954_ _13924_/A _13930_/X _13933_/A _13931_/Y VGND VGND VPWR VPWR _13954_/X sky130_fd_sc_hd__o22a_4
X_16742_ _22910_/A _16733_/Y _15991_/Y _23946_/Q VGND VGND VPWR VPWR _16742_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_6_43_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_87_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12905_ _12904_/X VGND VGND VPWR VPWR _25033_/D sky130_fd_sc_hd__inv_2
XFILLER_47_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16673_ _14754_/Y _16632_/A _16617_/X _16632_/A VGND VGND VPWR VPWR _24094_/D sky130_fd_sc_hd__a2bb2o_4
X_19461_ _19461_/A VGND VGND VPWR VPWR _19461_/Y sky130_fd_sc_hd__inv_2
X_13885_ _13885_/A VGND VGND VPWR VPWR _13886_/A sky130_fd_sc_hd__inv_2
X_18412_ _18412_/A _18452_/C VGND VGND VPWR VPWR _18440_/B sky130_fd_sc_hd__or2_4
X_12836_ _22396_/A VGND VGND VPWR VPWR _12836_/Y sky130_fd_sc_hd__inv_2
X_15624_ _15604_/A VGND VGND VPWR VPWR _15624_/X sky130_fd_sc_hd__buf_2
X_19392_ _15431_/X VGND VGND VPWR VPWR _19392_/X sky130_fd_sc_hd__buf_2
XFILLER_15_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23636__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15555_ _15553_/Y _15546_/X _15554_/X _15546_/X VGND VGND VPWR VPWR _24537_/D sky130_fd_sc_hd__a2bb2o_4
X_18343_ _18426_/C VGND VGND VPWR VPWR _18543_/A sky130_fd_sc_hd__buf_2
XANTENNA__15322__B _15531_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12767_ _12584_/Y _12762_/X VGND VGND VPWR VPWR _12767_/Y sky130_fd_sc_hd__nand2_4
XPHY_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14480_/X _14506_/B VGND VGND VPWR VPWR _14506_/X sky130_fd_sc_hd__or2_4
XPHY_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ _11707_/A _11718_/B VGND VGND VPWR VPWR _11719_/B sky130_fd_sc_hd__or2_4
X_18274_ _18279_/A _18278_/A _18202_/Y _18277_/B VGND VGND VPWR VPWR _18280_/B sky130_fd_sc_hd__or4_4
X_15486_ _12148_/Y _15475_/X _11558_/X _15475_/X VGND VGND VPWR VPWR _15486_/X sky130_fd_sc_hd__a2bb2o_4
X_12698_ _12636_/X VGND VGND VPWR VPWR _12716_/A sky130_fd_sc_hd__buf_2
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14437_ _14437_/A VGND VGND VPWR VPWR _14437_/X sky130_fd_sc_hd__buf_2
X_17225_ _11765_/A _11728_/X _11717_/A VGND VGND VPWR VPWR _18095_/B sky130_fd_sc_hd__and3_4
X_11649_ _13053_/A _11648_/X VGND VGND VPWR VPWR _11649_/Y sky130_fd_sc_hd__nand2_4
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17156_ _17086_/X _17134_/X _17156_/C VGND VGND VPWR VPWR _17156_/X sky130_fd_sc_hd__and3_4
X_14368_ _24768_/Q VGND VGND VPWR VPWR _14368_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16107_ _24332_/Q VGND VGND VPWR VPWR _16107_/Y sky130_fd_sc_hd__inv_2
X_13319_ _11735_/Y _13311_/X _13318_/X VGND VGND VPWR VPWR _13319_/X sky130_fd_sc_hd__and3_4
X_17087_ _17086_/X VGND VGND VPWR VPWR _17101_/A sky130_fd_sc_hd__buf_2
X_14299_ _24786_/Q VGND VGND VPWR VPWR _14299_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24495__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16038_ _11949_/Y _16038_/B _11512_/Y _16038_/D VGND VGND VPWR VPWR _16038_/X sky130_fd_sc_hd__or4_4
XFILLER_135_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24424__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_125_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_251_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17989_ _22272_/A _17987_/X _15788_/A _17987_/X VGND VGND VPWR VPWR _23920_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19728_ _11850_/A VGND VGND VPWR VPWR _19728_/X sky130_fd_sc_hd__buf_2
XFILLER_26_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21515__A _21224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19659_ _19646_/Y VGND VGND VPWR VPWR _19659_/X sky130_fd_sc_hd__buf_2
XFILLER_53_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15513__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22670_ _14860_/Y _21544_/X _14958_/Y _22312_/B VGND VGND VPWR VPWR _22670_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21621_ _17651_/A _21621_/B VGND VGND VPWR VPWR _21621_/X sky130_fd_sc_hd__or2_4
XANTENNA__25212__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21724__A2_N _21707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22340__B1 _11532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_63_0_HCLK clkbuf_8_63_0_HCLK/A VGND VGND VPWR VPWR _24361_/CLK sky130_fd_sc_hd__clkbuf_1
X_24340_ _24222_/CLK _24340_/D HRESETn VGND VGND VPWR VPWR _24340_/Q sky130_fd_sc_hd__dfrtp_4
X_21552_ _24796_/Q _16134_/X _21549_/X _21550_/X _21551_/X VGND VGND VPWR VPWR _21552_/X
+ sky130_fd_sc_hd__a2111o_4
X_20503_ _20502_/X VGND VGND VPWR VPWR _20503_/Y sky130_fd_sc_hd__inv_2
X_24271_ _24138_/CLK _16271_/X HRESETn VGND VGND VPWR VPWR _24271_/Q sky130_fd_sc_hd__dfrtp_4
X_21483_ _21350_/A _21481_/X _21482_/X VGND VGND VPWR VPWR _21483_/X sky130_fd_sc_hd__and3_4
XFILLER_105_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22025__A1_N _14223_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23222_ _23388_/CLK _23222_/D VGND VGND VPWR VPWR _19757_/A sky130_fd_sc_hd__dfxtp_4
X_20434_ _13503_/A _13503_/B _20433_/Y VGND VGND VPWR VPWR _20434_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__21446__A2 _20931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17159__B _17053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23153_ _23135_/CLK _19940_/X VGND VGND VPWR VPWR _23153_/Q sky130_fd_sc_hd__dfxtp_4
X_20365_ _14050_/Y _20344_/X _20358_/X _20364_/X VGND VGND VPWR VPWR _20365_/X sky130_fd_sc_hd__a211o_4
X_22104_ _20967_/A _22102_/X _22103_/X VGND VGND VPWR VPWR _22104_/X sky130_fd_sc_hd__and3_4
X_20296_ _20296_/A VGND VGND VPWR VPWR _20296_/X sky130_fd_sc_hd__buf_2
XFILLER_122_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24165__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23084_ _23085_/CLK _20120_/X VGND VGND VPWR VPWR _23084_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_115_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14884__B2 _22312_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22035_ _14012_/Y _14016_/X _23655_/Q _21088_/X VGND VGND VPWR VPWR _22039_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19272__B1 _19201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23986_ _23986_/CLK _17423_/X HRESETn VGND VGND VPWR VPWR _17253_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_113_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22937_ _22936_/X VGND VGND VPWR VPWR _22937_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13670_ _13408_/Y _13667_/X _13632_/X _13667_/X VGND VGND VPWR VPWR _24929_/D sky130_fd_sc_hd__a2bb2o_4
X_22868_ _13512_/C _22285_/X _23753_/Q _22531_/X VGND VGND VPWR VPWR _22868_/Y sky130_fd_sc_hd__a22oi_4
X_12621_ _25059_/Q _12619_/Y _12701_/A _24522_/Q VGND VGND VPWR VPWR _12622_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24607_ _24182_/CLK _24607_/D HRESETn VGND VGND VPWR VPWR _24607_/Q sky130_fd_sc_hd__dfrtp_4
X_21819_ _20979_/A _19602_/Y VGND VGND VPWR VPWR _21820_/C sky130_fd_sc_hd__or2_4
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22799_ _22799_/A VGND VGND VPWR VPWR _22799_/Y sky130_fd_sc_hd__inv_2
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15340_ _15353_/A VGND VGND VPWR VPWR _15340_/X sky130_fd_sc_hd__buf_2
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12552_ _12543_/X _12545_/X _12552_/C _12552_/D VGND VGND VPWR VPWR _12552_/X sky130_fd_sc_hd__or4_4
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24538_ _23486_/CLK _24538_/D HRESETn VGND VGND VPWR VPWR _19825_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22882__A1 _24249_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22256__A _22256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11503_ _11503_/A VGND VGND VPWR VPWR _21298_/B sky130_fd_sc_hd__buf_2
XFILLER_40_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15271_ _15271_/A _17197_/B VGND VGND VPWR VPWR _15285_/A sky130_fd_sc_hd__nor2_4
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12483_ _12460_/A _12478_/X _12483_/C VGND VGND VPWR VPWR _12483_/X sky130_fd_sc_hd__and3_4
X_24469_ _24488_/CLK _24469_/D HRESETn VGND VGND VPWR VPWR _12349_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16686__A2_N _16685_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16254__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24935__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17010_ _24049_/Q VGND VGND VPWR VPWR _17076_/A sky130_fd_sc_hd__inv_2
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14222_ _20332_/A _14201_/X _14221_/X _14201_/X VGND VGND VPWR VPWR _14222_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21437__A2 _20931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14153_ _12051_/A _12045_/X VGND VGND VPWR VPWR _14153_/X sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_5_27_0_HCLK_A clkbuf_5_27_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13104_ _13182_/A _13104_/B VGND VGND VPWR VPWR _13104_/X sky130_fd_sc_hd__or2_4
XFILLER_125_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14084_ _14079_/A VGND VGND VPWR VPWR _14084_/X sky130_fd_sc_hd__buf_2
X_18961_ _17935_/B VGND VGND VPWR VPWR _18961_/Y sky130_fd_sc_hd__inv_2
X_13035_ _13031_/X _13034_/X _11749_/X VGND VGND VPWR VPWR _13035_/X sky130_fd_sc_hd__o21a_4
X_17912_ _17944_/A _23464_/Q VGND VGND VPWR VPWR _17912_/X sky130_fd_sc_hd__or2_4
X_18892_ _18890_/Y _18891_/X _18823_/X _18891_/X VGND VGND VPWR VPWR _18892_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16077__B1 _15772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15419__A3 _15416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12350__A2 _12349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17843_ _15730_/X _17824_/X _17842_/X _23931_/Q _17765_/X VGND VGND VPWR VPWR _17843_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_66_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12323__A2_N _20808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23888__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17774_ _17887_/A _17774_/B VGND VGND VPWR VPWR _17774_/X sky130_fd_sc_hd__or2_4
X_14986_ _14986_/A VGND VGND VPWR VPWR _14986_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23817__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19513_ _23309_/Q VGND VGND VPWR VPWR _19513_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19551__A2_N _19546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16725_ _15965_/Y _22434_/A _15965_/Y _22434_/A VGND VGND VPWR VPWR _16725_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21335__A _21335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13937_ _13937_/A VGND VGND VPWR VPWR _13937_/X sky130_fd_sc_hd__buf_2
XFILLER_90_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22570__B1 _20777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19444_ _23333_/Q VGND VGND VPWR VPWR _21942_/B sky130_fd_sc_hd__inv_2
XFILLER_35_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13868_ _13868_/A VGND VGND VPWR VPWR _14352_/A sky130_fd_sc_hd__inv_2
X_16656_ _16655_/Y _16650_/X _15501_/X _16650_/X VGND VGND VPWR VPWR _24106_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11861__B2 _11830_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12819_ _21269_/A VGND VGND VPWR VPWR _12819_/Y sky130_fd_sc_hd__inv_2
X_15607_ _15604_/A VGND VGND VPWR VPWR _15607_/X sky130_fd_sc_hd__buf_2
XFILLER_37_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19375_ _13104_/B VGND VGND VPWR VPWR _19375_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21125__A1 _13357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13799_ scl_oen_o_S5 _13793_/X _13794_/Y _13798_/Y VGND VGND VPWR VPWR _13800_/B
+ sky130_fd_sc_hd__o22a_4
X_16587_ _16584_/A VGND VGND VPWR VPWR _16587_/X sky130_fd_sc_hd__buf_2
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18326_ _18167_/Y _18299_/X VGND VGND VPWR VPWR _18327_/B sky130_fd_sc_hd__or2_4
X_15538_ _15534_/Y _15537_/X RsRx_S0 _15537_/X VGND VGND VPWR VPWR _15538_/X sky130_fd_sc_hd__a2bb2o_4
X_15469_ _15368_/X _15461_/X _15468_/X _24575_/Q _15466_/X VGND VGND VPWR VPWR _15469_/X
+ sky130_fd_sc_hd__a32o_4
X_18257_ _18226_/A _18257_/B _18257_/C VGND VGND VPWR VPWR _23868_/D sky130_fd_sc_hd__and3_4
XFILLER_54_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16164__A _24310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24676__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17208_ _17208_/A VGND VGND VPWR VPWR _17208_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22625__A1 _22011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18188_ _16054_/A _18179_/Y _16116_/Y _23849_/Q VGND VGND VPWR VPWR _18190_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24605__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17139_ _17129_/A _17139_/B _17138_/X VGND VGND VPWR VPWR _24038_/D sky130_fd_sc_hd__and3_4
X_20150_ _23070_/Q VGND VGND VPWR VPWR _20150_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22389__B1 _24408_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20081_ _23099_/Q VGND VGND VPWR VPWR _20081_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17723__A _17716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23840_ _23840_/CLK _23840_/D HRESETn VGND VGND VPWR VPWR _23840_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21245__A _22564_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23771_ _23767_/CLK _20224_/X HRESETn VGND VGND VPWR VPWR _23771_/Q sky130_fd_sc_hd__dfrtp_4
X_20983_ _20961_/A _20983_/B VGND VGND VPWR VPWR _20983_/X sky130_fd_sc_hd__or2_4
XFILLER_53_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21364__A1 _22806_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16339__A _16339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22722_ _22943_/A _22721_/X VGND VGND VPWR VPWR _22722_/Y sky130_fd_sc_hd__nor2_4
XFILLER_81_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22653_ _12412_/C _22606_/X _24046_/Q _22652_/X VGND VGND VPWR VPWR _22659_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21604_ _17646_/A VGND VGND VPWR VPWR _21625_/A sky130_fd_sc_hd__buf_2
XFILLER_55_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22584_ _22584_/A VGND VGND VPWR VPWR _22585_/A sky130_fd_sc_hd__inv_2
X_24323_ _24071_/CLK _16128_/X HRESETn VGND VGND VPWR VPWR _20736_/A sky130_fd_sc_hd__dfrtp_4
X_21535_ _22146_/B _21533_/X _21256_/X _21534_/X VGND VGND VPWR VPWR _21535_/X sky130_fd_sc_hd__a211o_4
XFILLER_138_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24254_ _23767_/CLK _16303_/X HRESETn VGND VGND VPWR VPWR _16296_/A sky130_fd_sc_hd__dfrtp_4
X_21466_ _21469_/A _20086_/Y VGND VGND VPWR VPWR _21466_/X sky130_fd_sc_hd__or2_4
XANTENNA__24346__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_7_0_HCLK clkbuf_6_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_23205_ _24008_/CLK _23205_/D VGND VGND VPWR VPWR _13085_/B sky130_fd_sc_hd__dfxtp_4
X_20417_ _20414_/A _13517_/Y VGND VGND VPWR VPWR _20425_/A sky130_fd_sc_hd__or2_4
X_24185_ _24185_/CLK _16489_/X HRESETn VGND VGND VPWR VPWR _16488_/A sky130_fd_sc_hd__dfrtp_4
X_21397_ _21381_/X _21396_/X _21246_/X VGND VGND VPWR VPWR _21397_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__15649__A3 _15635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23136_ _25106_/CLK _19985_/X VGND VGND VPWR VPWR _23136_/Q sky130_fd_sc_hd__dfxtp_4
X_20348_ _20348_/A _20345_/A VGND VGND VPWR VPWR _20350_/B sky130_fd_sc_hd__nand2_4
XFILLER_107_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14857__B2 _24156_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15418__A _15418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11946__A _11507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23067_ _24013_/CLK _20550_/A VGND VGND VPWR VPWR _23067_/Q sky130_fd_sc_hd__dfxtp_4
X_20279_ _20279_/A _20279_/B _20278_/X VGND VGND VPWR VPWR _20279_/X sky130_fd_sc_hd__and3_4
X_22018_ _14916_/Y _22018_/B VGND VGND VPWR VPWR _22018_/X sky130_fd_sc_hd__and2_4
XFILLER_130_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23981__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14840_ _24699_/Q _14838_/Y _14839_/Y _14831_/A VGND VGND VPWR VPWR _14840_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23910__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14771_ _14770_/Y VGND VGND VPWR VPWR _15045_/A sky130_fd_sc_hd__buf_2
XANTENNA__25134__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11983_ _11983_/A VGND VGND VPWR VPWR _11983_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17559__B1 _16748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23969_ _23969_/CLK _17527_/X HRESETn VGND VGND VPWR VPWR _16693_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22552__B1 _16080_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13722_ _13722_/A VGND VGND VPWR VPWR _13722_/X sky130_fd_sc_hd__buf_2
X_16510_ _24176_/Q VGND VGND VPWR VPWR _16510_/Y sky130_fd_sc_hd__inv_2
X_17490_ _17490_/A _17490_/B VGND VGND VPWR VPWR _17491_/D sky130_fd_sc_hd__or2_4
XFILLER_95_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13653_ _13450_/Y _13649_/X _11590_/X _13652_/X VGND VGND VPWR VPWR _24938_/D sky130_fd_sc_hd__a2bb2o_4
X_16441_ _16441_/A VGND VGND VPWR VPWR _16441_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22304__B1 _24556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12604_ _12731_/A _24515_/Q _12731_/A _24515_/Q VGND VGND VPWR VPWR _12604_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16372_ _16364_/A VGND VGND VPWR VPWR _16372_/X sky130_fd_sc_hd__buf_2
X_19160_ _19153_/A VGND VGND VPWR VPWR _19160_/X sky130_fd_sc_hd__buf_2
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13584_ _13563_/X _13580_/X _13583_/Y _13576_/X _11673_/A VGND VGND VPWR VPWR _13584_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21602__B _21569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15323_ _11533_/X _15319_/Y _15320_/X _23026_/A _15325_/A VGND VGND VPWR VPWR _15323_/X
+ sky130_fd_sc_hd__a32o_4
X_18111_ _25137_/Q _18111_/B _18111_/C _12045_/X VGND VGND VPWR VPWR _18112_/A sky130_fd_sc_hd__or4_4
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12535_ _12456_/X _12535_/B _12534_/Y VGND VGND VPWR VPWR _25072_/D sky130_fd_sc_hd__and3_4
XFILLER_40_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19091_ _19091_/A VGND VGND VPWR VPWR _19091_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13621__A2_N _13620_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15254_ _15262_/A VGND VGND VPWR VPWR _15254_/X sky130_fd_sc_hd__buf_2
X_18042_ _23939_/Q VGND VGND VPWR VPWR _18043_/A sky130_fd_sc_hd__buf_2
X_12466_ _12413_/D _12466_/B VGND VGND VPWR VPWR _12467_/B sky130_fd_sc_hd__or2_4
XANTENNA__22607__B2 _22121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24087__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14205_ _14204_/Y _14200_/X _13665_/X _14202_/X VGND VGND VPWR VPWR _14205_/X sky130_fd_sc_hd__a2bb2o_4
X_15185_ _15184_/X VGND VGND VPWR VPWR _24664_/D sky130_fd_sc_hd__inv_2
XANTENNA__24016__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12397_ _12365_/X _12376_/X _12397_/C _12396_/X VGND VGND VPWR VPWR _12397_/X sky130_fd_sc_hd__or4_4
XANTENNA__16712__A _22202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14136_ _14126_/X _14135_/X _24991_/Q _14131_/X VGND VGND VPWR VPWR _14136_/X sky130_fd_sc_hd__o22a_4
X_19993_ _23133_/Q VGND VGND VPWR VPWR _19993_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14067_ _13764_/X _13742_/B _13742_/C _14066_/Y VGND VGND VPWR VPWR _14067_/X sky130_fd_sc_hd__and4_4
X_18944_ _18943_/X VGND VGND VPWR VPWR _18958_/A sky130_fd_sc_hd__buf_2
XANTENNA__14232__A _16373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13018_ _11753_/A _13018_/B _13017_/X VGND VGND VPWR VPWR _13018_/X sky130_fd_sc_hd__and3_4
XFILLER_80_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18875_ _18920_/A _19144_/B _18874_/X VGND VGND VPWR VPWR _18875_/X sky130_fd_sc_hd__or3_4
XFILLER_121_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17826_ _17861_/A _18792_/A VGND VGND VPWR VPWR _17826_/X sky130_fd_sc_hd__or2_4
XFILLER_67_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23651__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16470__B1 _16291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21065__A _21064_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17757_ _17928_/A _17757_/B VGND VGND VPWR VPWR _17757_/X sky130_fd_sc_hd__or2_4
XANTENNA__12087__B2 _24571_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14969_ _14969_/A VGND VGND VPWR VPWR _14969_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_5_13_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__22543__B1 _17558_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16708_ _23961_/Q VGND VGND VPWR VPWR _16708_/Y sky130_fd_sc_hd__inv_2
X_17688_ _17739_/A _17680_/X _17687_/X VGND VGND VPWR VPWR _17688_/X sky130_fd_sc_hd__or3_4
X_19427_ _13187_/B VGND VGND VPWR VPWR _19427_/Y sky130_fd_sc_hd__inv_2
X_16639_ _16632_/A VGND VGND VPWR VPWR _16639_/X sky130_fd_sc_hd__buf_2
XFILLER_23_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24857__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19358_ _19357_/Y _19355_/X _19221_/X _19355_/X VGND VGND VPWR VPWR _23363_/D sky130_fd_sc_hd__a2bb2o_4
X_18309_ _18212_/Y _18311_/B _18308_/Y VGND VGND VPWR VPWR _18309_/X sky130_fd_sc_hd__o21a_4
X_19289_ _19283_/Y VGND VGND VPWR VPWR _19289_/X sky130_fd_sc_hd__buf_2
X_21320_ _12534_/A _15456_/X _21319_/X VGND VGND VPWR VPWR _21320_/X sky130_fd_sc_hd__o21a_4
XFILLER_136_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13311__A _13073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_137_0_HCLK clkbuf_7_68_0_HCLK/X VGND VGND VPWR VPWR _23440_/CLK sky130_fd_sc_hd__clkbuf_1
X_21251_ _21251_/A _20826_/X VGND VGND VPWR VPWR _21251_/X sky130_fd_sc_hd__or2_4
XANTENNA__17718__A _17727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16622__A _16627_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22343__B _22281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16289__B1 _24258_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20202_ _23772_/Q VGND VGND VPWR VPWR _20202_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21182_ _20127_/Y _20827_/X VGND VGND VPWR VPWR _21182_/X sky130_fd_sc_hd__or2_4
XFILLER_137_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20133_ _23076_/Q VGND VGND VPWR VPWR _20133_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23739__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20064_ _23105_/Q VGND VGND VPWR VPWR _20064_/X sky130_fd_sc_hd__buf_2
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22997__C _22990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24941_ _24071_/CLK _24941_/D HRESETn VGND VGND VPWR VPWR _23036_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21585__A1 _11890_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24872_ _23676_/CLK _24872_/D HRESETn VGND VGND VPWR VPWR _20405_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15264__A1 _23766_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16461__B1 _16373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23823_ _23826_/CLK _23823_/D HRESETn VGND VGND VPWR VPWR _23823_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_72_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23754_ _24182_/CLK _23754_/D HRESETn VGND VGND VPWR VPWR _13540_/A sky130_fd_sc_hd__dfrtp_4
X_20966_ _20966_/A _20966_/B VGND VGND VPWR VPWR _20967_/C sky130_fd_sc_hd__or2_4
XFILLER_14_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22705_ _22597_/A _22704_/X VGND VGND VPWR VPWR _22705_/X sky130_fd_sc_hd__and2_4
XFILLER_96_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21703__A _21694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23685_ _23661_/CLK _23685_/D HRESETn VGND VGND VPWR VPWR _23685_/Q sky130_fd_sc_hd__dfstp_4
X_20897_ _20897_/A VGND VGND VPWR VPWR _20897_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24598__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22518__B _21979_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22636_ _22597_/A _22635_/X VGND VGND VPWR VPWR _22636_/X sky130_fd_sc_hd__and2_4
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24527__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19702__B2 _19701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16641__A1_N _14779_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_33_0_HCLK clkbuf_6_16_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_67_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22567_ _22681_/A _22564_/X _22566_/X VGND VGND VPWR VPWR _22567_/X sky130_fd_sc_hd__and3_4
X_12320_ _24494_/Q VGND VGND VPWR VPWR _12320_/Y sky130_fd_sc_hd__inv_2
X_24306_ _24308_/CLK _16175_/X HRESETn VGND VGND VPWR VPWR _24306_/Q sky130_fd_sc_hd__dfrtp_4
X_21518_ _21229_/A _21518_/B VGND VGND VPWR VPWR _21518_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_96_0_HCLK clkbuf_6_48_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_96_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__24180__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22498_ _15363_/Y _22497_/B VGND VGND VPWR VPWR _22498_/X sky130_fd_sc_hd__and2_4
XFILLER_120_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12251_ _25117_/Q _12250_/Y VGND VGND VPWR VPWR _12251_/X sky130_fd_sc_hd__or2_4
X_24237_ _24244_/CLK _24237_/D HRESETn VGND VGND VPWR VPWR _24237_/Q sky130_fd_sc_hd__dfrtp_4
X_21449_ _14043_/Y _14015_/A _24867_/Q _20844_/B VGND VGND VPWR VPWR _21449_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16656__A1_N _16655_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12182_ _12132_/Y _12127_/Y _12256_/B VGND VGND VPWR VPWR _12183_/B sky130_fd_sc_hd__or3_4
X_24168_ _24168_/CLK _16531_/X HRESETn VGND VGND VPWR VPWR _24168_/Q sky130_fd_sc_hd__dfrtp_4
X_23119_ _23401_/CLK _20030_/X VGND VGND VPWR VPWR _20029_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_123_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_16990_ _16990_/A _16990_/B _16987_/X _16989_/X VGND VGND VPWR VPWR _16991_/D sky130_fd_sc_hd__or4_4
XFILLER_1_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24099_ _24098_/CLK _16667_/X HRESETn VGND VGND VPWR VPWR _24099_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15941_ _15928_/X VGND VGND VPWR VPWR _15941_/X sky130_fd_sc_hd__buf_2
XFILLER_114_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18459__A _18459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18660_ _18659_/Y _18657_/X _15566_/X _18657_/X VGND VGND VPWR VPWR _18660_/X sky130_fd_sc_hd__a2bb2o_4
X_15872_ _24409_/Q VGND VGND VPWR VPWR _15872_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17611_ _17484_/Y _17587_/B _17528_/X _17609_/B VGND VGND VPWR VPWR _17611_/X sky130_fd_sc_hd__a211o_4
X_14823_ _24152_/Q VGND VGND VPWR VPWR _14823_/Y sky130_fd_sc_hd__inv_2
X_18591_ _16356_/Y _23825_/Q _16356_/Y _23825_/Q VGND VGND VPWR VPWR _18591_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22525__B1 _24411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17542_ _17481_/A _17545_/B VGND VGND VPWR VPWR _17542_/X sky130_fd_sc_hd__or2_4
X_11966_ _11965_/Y VGND VGND VPWR VPWR _11966_/X sky130_fd_sc_hd__buf_2
X_14754_ _14754_/A VGND VGND VPWR VPWR _14754_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16204__B1 _15894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22709__A _24310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13705_ _13697_/X _13704_/X _14090_/A _13682_/Y VGND VGND VPWR VPWR _13705_/X sky130_fd_sc_hd__o22a_4
X_14685_ _14059_/Y _14621_/X _14622_/X _14684_/X VGND VGND VPWR VPWR _14686_/A sky130_fd_sc_hd__o22a_4
X_17473_ _17461_/X _17457_/Y _17472_/X _21799_/A _17462_/Y VGND VGND VPWR VPWR _23975_/D
+ sky130_fd_sc_hd__a32o_4
X_11897_ _13370_/A _11896_/Y _13370_/A _11896_/Y VGND VGND VPWR VPWR _11902_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18194__A _18468_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24950__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19212_ _13611_/X _16127_/A VGND VGND VPWR VPWR _19212_/Y sky130_fd_sc_hd__nor2_4
X_13636_ _13634_/Y _13631_/X _13635_/X _13631_/X VGND VGND VPWR VPWR _24944_/D sky130_fd_sc_hd__a2bb2o_4
X_16424_ _16423_/Y _16421_/X _16259_/X _16421_/X VGND VGND VPWR VPWR _16424_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15611__A _16624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22828__A1 _17482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24268__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16609__A1_N _16608_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19143_ _17697_/B VGND VGND VPWR VPWR _19143_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13567_ _13567_/A _13567_/B VGND VGND VPWR VPWR _13568_/B sky130_fd_sc_hd__or2_4
X_16355_ _16354_/Y _16352_/X _16093_/X _16352_/X VGND VGND VPWR VPWR _16355_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17704__B1 _15712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18922__A _18935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14227__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12518_ _12328_/Y _12515_/B VGND VGND VPWR VPWR _12519_/C sky130_fd_sc_hd__nand2_4
X_15306_ _11950_/X _15304_/X HADDR[21] _15304_/X VGND VGND VPWR VPWR _15306_/X sky130_fd_sc_hd__a2bb2o_4
X_16286_ _16262_/A VGND VGND VPWR VPWR _16286_/X sky130_fd_sc_hd__buf_2
X_19074_ _19073_/Y _19071_/X _18938_/X _19071_/X VGND VGND VPWR VPWR _23464_/D sky130_fd_sc_hd__a2bb2o_4
X_13498_ _13498_/A VGND VGND VPWR VPWR _13498_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22444__A _24107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18025_ _18020_/X _18061_/B _18022_/X _18025_/D VGND VGND VPWR VPWR _18025_/X sky130_fd_sc_hd__and4_4
XFILLER_117_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12449_ _12451_/B VGND VGND VPWR VPWR _12449_/Y sky130_fd_sc_hd__inv_2
X_15237_ _13777_/X _15237_/B _13790_/X _14068_/X VGND VGND VPWR VPWR _15237_/X sky130_fd_sc_hd__or4_4
XANTENNA__21264__B1 _24547_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15168_ _14941_/Y _15159_/X VGND VGND VPWR VPWR _15168_/X sky130_fd_sc_hd__or2_4
X_14119_ _14119_/A VGND VGND VPWR VPWR _14120_/B sky130_fd_sc_hd__inv_2
XFILLER_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15099_ _15099_/A VGND VGND VPWR VPWR _15159_/A sky130_fd_sc_hd__inv_2
X_19976_ _21777_/B _19970_/X _19448_/A _19975_/X VGND VGND VPWR VPWR _19976_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20899__A _21109_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23832__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24804__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18927_ _18935_/A VGND VGND VPWR VPWR _18927_/X sky130_fd_sc_hd__buf_2
XANTENNA__25056__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24867__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18858_ _23540_/Q VGND VGND VPWR VPWR _18858_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17809_ _17879_/A _17809_/B _17809_/C VGND VGND VPWR VPWR _17815_/B sky130_fd_sc_hd__and3_4
X_18789_ _23564_/Q VGND VGND VPWR VPWR _18789_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21319__A1 _17615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22516__B1 _24561_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20820_ _20819_/X VGND VGND VPWR VPWR _20820_/X sky130_fd_sc_hd__buf_2
XFILLER_36_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20751_ _11501_/X VGND VGND VPWR VPWR _20751_/X sky130_fd_sc_hd__buf_2
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24691__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16617__A _16216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23470_ _24733_/CLK _23470_/D VGND VGND VPWR VPWR _23470_/Q sky130_fd_sc_hd__dfxtp_4
X_20682_ _20556_/X _20681_/X _24188_/Q _20602_/X VGND VGND VPWR VPWR _23757_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24620__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22421_ _24516_/Q _20799_/X _20801_/X _22420_/X VGND VGND VPWR VPWR _22421_/X sky130_fd_sc_hd__a211o_4
XFILLER_91_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25140_ _25141_/CLK _25140_/D HRESETn VGND VGND VPWR VPWR _25140_/Q sky130_fd_sc_hd__dfrtp_4
X_22352_ _24336_/Q _22350_/X _22351_/X VGND VGND VPWR VPWR _22352_/X sky130_fd_sc_hd__o21a_4
XFILLER_104_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21303_ _13376_/Y _20751_/X _11930_/Y _21083_/X VGND VGND VPWR VPWR _21303_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11991__B1 _11604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25071_ _25097_/CLK _12537_/X HRESETn VGND VGND VPWR VPWR _21104_/A sky130_fd_sc_hd__dfrtp_4
X_22283_ _20927_/X _22278_/X _22280_/X _22282_/X VGND VGND VPWR VPWR _22284_/B sky130_fd_sc_hd__o22a_4
XFILLER_117_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24022_ _23664_/CLK _17193_/X HRESETn VGND VGND VPWR VPWR _24022_/Q sky130_fd_sc_hd__dfstp_4
X_21234_ _21234_/A VGND VGND VPWR VPWR _21235_/A sky130_fd_sc_hd__buf_2
XFILLER_89_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11496__A _11496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21165_ _21153_/A VGND VGND VPWR VPWR _21935_/A sky130_fd_sc_hd__buf_2
XANTENNA__16277__A3 _16100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20116_ _17979_/X _21795_/B VGND VGND VPWR VPWR _20116_/X sky130_fd_sc_hd__or2_4
X_21096_ _21275_/A VGND VGND VPWR VPWR _21719_/A sky130_fd_sc_hd__buf_2
XANTENNA__20602__A _20651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20047_ _20047_/A VGND VGND VPWR VPWR _21342_/B sky130_fd_sc_hd__inv_2
XFILLER_59_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24924_ _24879_/CLK _24924_/D HRESETn VGND VGND VPWR VPWR _20201_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_115_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24855_ _23657_/CLK _24855_/D HRESETn VGND VGND VPWR VPWR _14096_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22507__B1 _20821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24779__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11820_ _11776_/B _11817_/B VGND VGND VPWR VPWR _11824_/A sky130_fd_sc_hd__and2_4
XANTENNA__13216__A _13092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13799__A1 scl_oen_o_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23806_ _23648_/CLK _23806_/D HRESETn VGND VGND VPWR VPWR _20705_/B sky130_fd_sc_hd__dfstp_4
X_24786_ _24776_/CLK _24786_/D HRESETn VGND VGND VPWR VPWR _24786_/Q sky130_fd_sc_hd__dfrtp_4
X_21998_ _16961_/A _21066_/B VGND VGND VPWR VPWR _22002_/B sky130_fd_sc_hd__and2_4
XANTENNA__24708__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11732_/A VGND VGND VPWR VPWR _11751_/X sky130_fd_sc_hd__buf_2
XPHY_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23737_ _24259_/CLK _23737_/D HRESETn VGND VGND VPWR VPWR _23737_/Q sky130_fd_sc_hd__dfrtp_4
X_20949_ _17642_/Y VGND VGND VPWR VPWR _21626_/A sky130_fd_sc_hd__buf_2
XANTENNA__21730__A1 _21562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15431__A HWDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _14469_/X VGND VGND VPWR VPWR _14471_/A sky130_fd_sc_hd__inv_2
XANTENNA__14748__B1 _15087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11682_/A _11682_/B _11682_/C _11681_/X VGND VGND VPWR VPWR _11694_/C sky130_fd_sc_hd__or4_4
XANTENNA__16580__A1_N _14850_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24361__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23668_ _23668_/CLK _20352_/Y HRESETn VGND VGND VPWR VPWR _20348_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _24926_/Q VGND VGND VPWR VPWR _13421_/Y sky130_fd_sc_hd__inv_2
XPHY_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22619_ _22691_/A _22619_/B _22619_/C VGND VGND VPWR VPWR _22661_/A sky130_fd_sc_hd__and3_4
XFILLER_70_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22286__A2 _22173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14047__A _14047_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23599_ _23992_/CLK _18688_/X VGND VGND VPWR VPWR _13300_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_31_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16140_ _24319_/Q VGND VGND VPWR VPWR _16140_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13352_ _13350_/Y _13351_/X _11636_/X _13351_/X VGND VGND VPWR VPWR _24989_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21494__B1 _23913_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12303_ _25081_/Q VGND VGND VPWR VPWR _12508_/A sky130_fd_sc_hd__inv_2
XANTENNA__11982__B1 _11981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16071_ _16071_/A VGND VGND VPWR VPWR _16071_/X sky130_fd_sc_hd__buf_2
XFILLER_6_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13283_ _13219_/A _13283_/B VGND VGND VPWR VPWR _13283_/X sky130_fd_sc_hd__or2_4
XFILLER_127_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15022_ _15022_/A _15021_/X VGND VGND VPWR VPWR _15025_/B sky130_fd_sc_hd__or2_4
Xclkbuf_8_120_0_HCLK clkbuf_7_60_0_HCLK/X VGND VGND VPWR VPWR _23852_/CLK sky130_fd_sc_hd__clkbuf_1
X_12234_ _12227_/X _12234_/B _12233_/X VGND VGND VPWR VPWR _12234_/X sky130_fd_sc_hd__and3_4
XFILLER_120_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_183_0_HCLK clkbuf_7_91_0_HCLK/X VGND VGND VPWR VPWR _24478_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_135_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22994__B1 _22530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19830_ _23193_/Q VGND VGND VPWR VPWR _19830_/Y sky130_fd_sc_hd__inv_2
X_12165_ _12418_/C VGND VGND VPWR VPWR _12165_/X sky130_fd_sc_hd__buf_2
XFILLER_122_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16673__B1 _16617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19761_ _22095_/B _19760_/X _19711_/X _19760_/X VGND VGND VPWR VPWR _23222_/D sky130_fd_sc_hd__a2bb2o_4
X_12096_ _25121_/Q _24564_/Q _12094_/Y _12095_/Y VGND VGND VPWR VPWR _12096_/X sky130_fd_sc_hd__o22a_4
X_16973_ _24045_/Q VGND VGND VPWR VPWR _17042_/A sky130_fd_sc_hd__inv_2
X_18712_ _18711_/X VGND VGND VPWR VPWR _18712_/X sky130_fd_sc_hd__buf_2
X_15924_ _15918_/Y _15923_/X _15828_/X _15923_/X VGND VGND VPWR VPWR _15924_/X sky130_fd_sc_hd__a2bb2o_4
X_19692_ _19691_/Y _19689_/X _19600_/X _19689_/X VGND VGND VPWR VPWR _23245_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18643_ _14540_/X _19862_/B _19883_/C VGND VGND VPWR VPWR _18644_/A sky130_fd_sc_hd__or3_4
X_15855_ HWDATA[21] VGND VGND VPWR VPWR _15855_/X sky130_fd_sc_hd__buf_2
XFILLER_92_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13126__A _13073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14806_ _14703_/X _24150_/Q _14703_/X _24150_/Q VGND VGND VPWR VPWR _14806_/X sky130_fd_sc_hd__a2bb2o_4
X_18574_ _16366_/A _23821_/Q _16366_/Y _18536_/A VGND VGND VPWR VPWR _18574_/X sky130_fd_sc_hd__o22a_4
X_15786_ _15781_/X _15582_/A _16100_/A _24440_/Q _15746_/A VGND VGND VPWR VPWR _24440_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_52_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24449__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12998_ _12793_/Y _12915_/C VGND VGND VPWR VPWR _13008_/B sky130_fd_sc_hd__or2_4
XANTENNA__22439__A _16351_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18636__B _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17525_ _16693_/A _17524_/Y VGND VGND VPWR VPWR _17525_/X sky130_fd_sc_hd__or2_4
XFILLER_73_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14737_ _14737_/A VGND VGND VPWR VPWR _14737_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11949_ _11949_/A VGND VGND VPWR VPWR _11949_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16728__B2 _17481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21721__B2 _20757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17456_ _17455_/Y _17453_/A _21799_/A _17452_/A VGND VGND VPWR VPWR _17457_/B sky130_fd_sc_hd__o22a_4
XFILLER_60_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14668_ _14640_/X _14667_/X _14050_/A _14647_/X VGND VGND VPWR VPWR _14668_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16407_ _16406_/Y _16402_/X _16246_/X _16402_/X VGND VGND VPWR VPWR _16407_/X sky130_fd_sc_hd__a2bb2o_4
X_13619_ _16305_/A VGND VGND VPWR VPWR _13619_/X sky130_fd_sc_hd__buf_2
X_17387_ _17266_/Y _17386_/X VGND VGND VPWR VPWR _17388_/C sky130_fd_sc_hd__nand2_4
XANTENNA__24031__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14599_ _24733_/Q VGND VGND VPWR VPWR _19123_/B sky130_fd_sc_hd__buf_2
X_19126_ _19122_/Y _19125_/X _19059_/X _19125_/X VGND VGND VPWR VPWR _23446_/D sky130_fd_sc_hd__a2bb2o_4
X_16338_ _24241_/Q VGND VGND VPWR VPWR _16338_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19057_ _18874_/X _19100_/B VGND VGND VPWR VPWR _19071_/A sky130_fd_sc_hd__nor2_4
X_16269_ _16234_/A VGND VGND VPWR VPWR _16269_/X sky130_fd_sc_hd__buf_2
XANTENNA__16172__A _16172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18008_ _18007_/Y VGND VGND VPWR VPWR _18008_/X sky130_fd_sc_hd__buf_2
XFILLER_133_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22378__A1_N _12495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22985__B1 _22840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19850__B1 _19825_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15467__A1 _15368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16664__B1 _16455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21518__A _21229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19959_ _23145_/Q VGND VGND VPWR VPWR _19959_/Y sky130_fd_sc_hd__inv_2
X_22970_ _22335_/A _22969_/X _22835_/X _11496_/A _22840_/X VGND VGND VPWR VPWR _22970_/X
+ sky130_fd_sc_hd__a32o_4
X_21921_ _20975_/A _21919_/X _21920_/X VGND VGND VPWR VPWR _21921_/X sky130_fd_sc_hd__and3_4
XANTENNA__24872__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13036__A _13011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24640_ _23762_/CLK _15261_/X HRESETn VGND VGND VPWR VPWR _24640_/Q sky130_fd_sc_hd__dfrtp_4
X_21852_ _21034_/Y VGND VGND VPWR VPWR _22629_/A sky130_fd_sc_hd__buf_2
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20803_ _24500_/Q _20826_/A _20739_/B _15642_/X VGND VGND VPWR VPWR _20803_/X sky130_fd_sc_hd__o22a_4
XFILLER_93_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24571_ _24488_/CLK _24571_/D HRESETn VGND VGND VPWR VPWR _24571_/Q sky130_fd_sc_hd__dfrtp_4
X_21783_ _21779_/X _21782_/X _14523_/A VGND VGND VPWR VPWR _21783_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__24119__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13650__B1 _11581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16719__B2 _23947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12875__A _22258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23522_ _23563_/CLK _18911_/X VGND VGND VPWR VPWR _17868_/B sky130_fd_sc_hd__dfxtp_4
X_20734_ sda_oen_o_S5 _24624_/Q _20729_/A _15234_/X _20733_/Y VGND VGND VPWR VPWR
+ _20734_/X sky130_fd_sc_hd__a32o_4
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23453_ _23469_/CLK _23453_/D VGND VGND VPWR VPWR _17712_/B sky130_fd_sc_hd__dfxtp_4
X_20665_ _20663_/Y _20660_/Y _20664_/X VGND VGND VPWR VPWR _20665_/X sky130_fd_sc_hd__o21a_4
XFILLER_50_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22404_ _22263_/X _22404_/B VGND VGND VPWR VPWR _22404_/Y sky130_fd_sc_hd__nor2_4
X_23384_ _23385_/CLK _19299_/X VGND VGND VPWR VPWR _19298_/A sky130_fd_sc_hd__dfxtp_4
X_20596_ _16532_/Y _20574_/X _20583_/X _20595_/X VGND VGND VPWR VPWR _20597_/A sky130_fd_sc_hd__o22a_4
XFILLER_104_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25123_ _25123_/CLK _12234_/X HRESETn VGND VGND VPWR VPWR _12172_/A sky130_fd_sc_hd__dfrtp_4
X_22335_ _22335_/A VGND VGND VPWR VPWR _22574_/B sky130_fd_sc_hd__buf_2
XFILLER_87_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16082__A _24340_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23754__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25054_ _24521_/CLK _12718_/X HRESETn VGND VGND VPWR VPWR _25054_/Q sky130_fd_sc_hd__dfrtp_4
X_22266_ _22264_/X _22265_/X _14831_/Y _16305_/X VGND VGND VPWR VPWR _22266_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11938__B _21300_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22812__A _22811_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22976__B1 _24575_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24005_ _24005_/CLK _17354_/X HRESETn VGND VGND VPWR VPWR _17352_/A sky130_fd_sc_hd__dfrtp_4
X_21217_ _21212_/X _21216_/X _14524_/D VGND VGND VPWR VPWR _21217_/X sky130_fd_sc_hd__o21a_4
XFILLER_104_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22197_ _22197_/A VGND VGND VPWR VPWR _22197_/X sky130_fd_sc_hd__buf_2
XANTENNA__14951__A1_N _14950_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17998__A3 _15704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21148_ _21144_/X _21147_/X _17639_/X VGND VGND VPWR VPWR _21148_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22728__B1 _16068_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15426__A _20861_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13970_ _13937_/X _13969_/X _14259_/A _13963_/X VGND VGND VPWR VPWR _13970_/Y sky130_fd_sc_hd__a22oi_4
X_21079_ _20852_/A _21079_/B VGND VGND VPWR VPWR _21079_/X sky130_fd_sc_hd__or2_4
XANTENNA__16670__A3 _15706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16407__B1 _16246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23065__D scl_oen_o_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12921_ _12921_/A _12921_/B _12920_/X VGND VGND VPWR VPWR _12921_/X sky130_fd_sc_hd__and3_4
XFILLER_111_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24907_ _24904_/CLK _13904_/X HRESETn VGND VGND VPWR VPWR _24907_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15640_ _15639_/X VGND VGND VPWR VPWR _22218_/C sky130_fd_sc_hd__buf_2
XFILLER_74_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12852_ _12788_/Y _24455_/Q _12854_/A _12851_/Y VGND VGND VPWR VPWR _12856_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24838_ _24851_/CLK _14152_/X HRESETn VGND VGND VPWR VPWR _24838_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24542__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22259__A _22259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11803_ _11799_/Y _11803_/B _11803_/C VGND VGND VPWR VPWR _11804_/A sky130_fd_sc_hd__or3_4
XFILLER_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12783_ _12775_/X _12783_/B _12780_/X _12782_/X VGND VGND VPWR VPWR _12783_/X sky130_fd_sc_hd__or4_4
X_15571_ _22884_/B VGND VGND VPWR VPWR _15572_/A sky130_fd_sc_hd__buf_2
XFILLER_92_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24769_ _24769_/CLK _24769_/D HRESETn VGND VGND VPWR VPWR _24769_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17310_/A VGND VGND VPWR VPWR _17312_/C sky130_fd_sc_hd__inv_2
XPHY_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11734_ _23897_/Q VGND VGND VPWR VPWR _11734_/Y sky130_fd_sc_hd__inv_2
X_14522_ _14440_/X VGND VGND VPWR VPWR _14523_/A sky130_fd_sc_hd__buf_2
XFILLER_109_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18290_ _18262_/A VGND VGND VPWR VPWR _18290_/X sky130_fd_sc_hd__buf_2
XPHY_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _11547_/Y _17306_/A _11547_/Y _17306_/A VGND VGND VPWR VPWR _17241_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _11665_/A VGND VGND VPWR VPWR _22319_/A sky130_fd_sc_hd__inv_2
X_14453_ _14524_/B _14452_/X _14524_/B _14452_/X VGND VGND VPWR VPWR _14453_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15394__B1 _15393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ _15807_/A VGND VGND VPWR VPWR _15712_/A sky130_fd_sc_hd__inv_2
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14384_ _13432_/Y _14402_/B VGND VGND VPWR VPWR _14384_/X sky130_fd_sc_hd__or2_4
X_17172_ _20348_/A _20345_/A VGND VGND VPWR VPWR _17173_/B sky130_fd_sc_hd__or2_4
XANTENNA__22177__A2_N _22857_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11596_ _25201_/Q VGND VGND VPWR VPWR _11596_/Y sky130_fd_sc_hd__inv_2
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13335_ _13334_/X VGND VGND VPWR VPWR _13335_/X sky130_fd_sc_hd__buf_2
X_16123_ _16123_/A VGND VGND VPWR VPWR _21097_/A sky130_fd_sc_hd__inv_2
X_13266_ _13202_/A _13266_/B VGND VGND VPWR VPWR _13267_/C sky130_fd_sc_hd__or2_4
X_16054_ _16054_/A VGND VGND VPWR VPWR _16054_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12217_ _12079_/X _12216_/X _12195_/X VGND VGND VPWR VPWR _12217_/Y sky130_fd_sc_hd__a21oi_4
X_15005_ _14868_/B _15014_/B VGND VGND VPWR VPWR _15006_/A sky130_fd_sc_hd__or2_4
XANTENNA__18635__A1 _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13197_ _13261_/A _13197_/B VGND VGND VPWR VPWR _13197_/X sky130_fd_sc_hd__or2_4
XFILLER_69_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19813_ _19813_/A VGND VGND VPWR VPWR _19831_/A sky130_fd_sc_hd__inv_2
XFILLER_29_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16646__B1 HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12148_ _24567_/Q VGND VGND VPWR VPWR _12148_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19744_ _21824_/B _19738_/X _19717_/X _19743_/X VGND VGND VPWR VPWR _19744_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12079_ _12078_/Y VGND VGND VPWR VPWR _12079_/X sky130_fd_sc_hd__buf_2
X_16956_ _16952_/B _16955_/X _16951_/C VGND VGND VPWR VPWR _24060_/D sky130_fd_sc_hd__and3_4
XFILLER_110_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15907_ _15906_/Y _15826_/X _15709_/X _15826_/X VGND VGND VPWR VPWR _24396_/D sky130_fd_sc_hd__a2bb2o_4
X_19675_ _23251_/Q VGND VGND VPWR VPWR _19675_/Y sky130_fd_sc_hd__inv_2
X_16887_ _16887_/A VGND VGND VPWR VPWR _16888_/B sky130_fd_sc_hd__inv_2
XFILLER_37_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20896__B _20868_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18626_ _18607_/X _18621_/X _23809_/Q _23810_/Q _18624_/X VGND VGND VPWR VPWR _18626_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17551__A _17497_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15838_ _15836_/Y _15834_/X _15837_/X _15834_/X VGND VGND VPWR VPWR _15838_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24283__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22169__A _22952_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18557_ _18551_/A _18551_/B VGND VGND VPWR VPWR _18558_/C sky130_fd_sc_hd__nand2_4
XFILLER_64_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12435__A1 _12401_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15769_ _12790_/Y _15768_/X _15350_/X _15768_/X VGND VGND VPWR VPWR _15769_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24212__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17508_ _23012_/A _17508_/B VGND VGND VPWR VPWR _17509_/C sky130_fd_sc_hd__nand2_4
XFILLER_75_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18488_ _18488_/A _18488_/B VGND VGND VPWR VPWR _18491_/B sky130_fd_sc_hd__or2_4
XFILLER_75_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17439_ _17264_/Y _17434_/X VGND VGND VPWR VPWR _17440_/B sky130_fd_sc_hd__nand2_4
XFILLER_123_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20450_ _20447_/Y _20442_/Y _20453_/B VGND VGND VPWR VPWR _20450_/X sky130_fd_sc_hd__o21a_4
XFILLER_88_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19109_ _16545_/X VGND VGND VPWR VPWR _19109_/X sky130_fd_sc_hd__buf_2
X_20381_ _23675_/Q _17179_/B VGND VGND VPWR VPWR _20381_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22670__A2 _21544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22120_ _22438_/A _22120_/B VGND VGND VPWR VPWR _22120_/X sky130_fd_sc_hd__and2_4
XFILLER_118_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25071__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22632__A _21848_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22051_ _21308_/X _22028_/X _22040_/X _22050_/X VGND VGND VPWR VPWR _22051_/X sky130_fd_sc_hd__a211o_4
XANTENNA__25000__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21002_ _21006_/A _21002_/B VGND VGND VPWR VPWR _21003_/C sky130_fd_sc_hd__or2_4
XFILLER_102_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16637__B1 _24116_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22973__A3 _22459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_23_0_HCLK clkbuf_8_23_0_HCLK/A VGND VGND VPWR VPWR _24757_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_101_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_86_0_HCLK clkbuf_8_87_0_HCLK/A VGND VGND VPWR VPWR _24897_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22953_ _24318_/Q _22953_/B VGND VGND VPWR VPWR _22953_/X sky130_fd_sc_hd__and2_4
X_21904_ _14050_/Y _20818_/A _14639_/A _20832_/A VGND VGND VPWR VPWR _21905_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22884_ _22884_/A _22884_/B VGND VGND VPWR VPWR _22884_/X sky130_fd_sc_hd__and2_4
XFILLER_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21835_ _22105_/A _21834_/X _23941_/Q VGND VGND VPWR VPWR _21835_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_43_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24623_ _24623_/CLK _24623_/D HRESETn VGND VGND VPWR VPWR _11505_/A sky130_fd_sc_hd__dfrtp_4
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24554_ _24566_/CLK _24554_/D HRESETn VGND VGND VPWR VPWR _24554_/Q sky130_fd_sc_hd__dfrtp_4
X_21766_ _21762_/X _21766_/B VGND VGND VPWR VPWR _21766_/X sky130_fd_sc_hd__or2_4
XFILLER_19_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17000__A2_N _24040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20717_ _20717_/A _23615_/Q VGND VGND VPWR VPWR _20717_/X sky130_fd_sc_hd__and2_4
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23505_ _23511_/CLK _23505_/D VGND VGND VPWR VPWR _17903_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24485_ _24488_/CLK _24485_/D HRESETn VGND VGND VPWR VPWR _22591_/A sky130_fd_sc_hd__dfrtp_4
X_21697_ _21700_/A _23394_/Q _13403_/A _19273_/Y VGND VGND VPWR VPWR _21697_/X sky130_fd_sc_hd__o22a_4
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21449__B1 _24867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23935__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23436_ _25067_/CLK _19154_/X VGND VGND VPWR VPWR _23436_/Q sky130_fd_sc_hd__dfxtp_4
X_20648_ _23748_/Q VGND VGND VPWR VPWR _20648_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21430__B _20818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25159__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14718__A2_N _24093_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23367_ _24998_/CLK _19346_/X VGND VGND VPWR VPWR _13305_/B sky130_fd_sc_hd__dfxtp_4
X_20579_ _13533_/B VGND VGND VPWR VPWR _20579_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17015__A2_N _17022_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13120_ _13078_/A VGND VGND VPWR VPWR _13120_/X sky130_fd_sc_hd__buf_2
X_22318_ _13655_/Y _20911_/X VGND VGND VPWR VPWR _22318_/X sky130_fd_sc_hd__and2_4
X_25106_ _25106_/CLK _25106_/D HRESETn VGND VGND VPWR VPWR _25106_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23298_ _23112_/CLK _23298_/D VGND VGND VPWR VPWR _19543_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_124_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22949__B1 _16050_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13051_ _13047_/X _13050_/X _11749_/X VGND VGND VPWR VPWR _13051_/X sky130_fd_sc_hd__o21a_4
X_25037_ _25044_/CLK _12773_/Y HRESETn VGND VGND VPWR VPWR _12562_/A sky130_fd_sc_hd__dfrtp_4
X_22249_ _22249_/A VGND VGND VPWR VPWR _22999_/B sky130_fd_sc_hd__buf_2
XFILLER_121_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22413__A2 _21882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22208__A1_N _11913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12002_ _11990_/A VGND VGND VPWR VPWR _12002_/X sky130_fd_sc_hd__buf_2
XFILLER_78_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19290__B2 _19289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24794__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16810_ _16791_/X _16796_/X _16804_/X _16810_/D VGND VGND VPWR VPWR _16811_/B sky130_fd_sc_hd__or4_4
X_17790_ _17918_/A VGND VGND VPWR VPWR _17929_/A sky130_fd_sc_hd__buf_2
XFILLER_66_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24723__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22177__B2 _16134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16741_ _15925_/Y _22979_/A _15925_/Y _22979_/A VGND VGND VPWR VPWR _16744_/B sky130_fd_sc_hd__a2bb2o_4
X_13953_ _13936_/A VGND VGND VPWR VPWR _13959_/A sky130_fd_sc_hd__buf_2
XFILLER_59_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12904_ _12899_/C _12894_/B _12896_/X _12900_/Y VGND VGND VPWR VPWR _12904_/X sky130_fd_sc_hd__a211o_4
X_19460_ _19457_/Y _19458_/X _19459_/X _19458_/X VGND VGND VPWR VPWR _23329_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17371__A _17303_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16672_ _14747_/Y _16666_/X _16671_/X _16666_/X VGND VGND VPWR VPWR _24095_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13884_ _13905_/A VGND VGND VPWR VPWR _13884_/X sky130_fd_sc_hd__buf_2
XFILLER_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18411_ _23843_/Q VGND VGND VPWR VPWR _18440_/A sky130_fd_sc_hd__inv_2
X_15623_ _12582_/Y _15621_/X _15511_/X _15621_/X VGND VGND VPWR VPWR _24511_/D sky130_fd_sc_hd__a2bb2o_4
X_12835_ _12825_/X _12828_/X _12835_/C _12835_/D VGND VGND VPWR VPWR _12835_/X sky130_fd_sc_hd__or4_4
X_19391_ _19391_/A VGND VGND VPWR VPWR _19391_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18342_ _23819_/Q VGND VGND VPWR VPWR _18426_/C sky130_fd_sc_hd__inv_2
X_15554_ _19452_/A VGND VGND VPWR VPWR _15554_/X sky130_fd_sc_hd__buf_2
X_12766_ _12766_/A _12766_/B _12755_/X VGND VGND VPWR VPWR _12766_/X sky130_fd_sc_hd__and3_4
XPHY_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18553__B1 _18449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _14502_/Y _14480_/X _14504_/Y VGND VGND VPWR VPWR _14505_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21621__A _17651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11717_ _11717_/A VGND VGND VPWR VPWR _21188_/A sky130_fd_sc_hd__buf_2
X_18273_ _18203_/Y _18273_/B VGND VGND VPWR VPWR _18277_/B sky130_fd_sc_hd__or2_4
XANTENNA__15367__B1 _11581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _12696_/X VGND VGND VPWR VPWR _25059_/D sky130_fd_sc_hd__inv_2
X_15485_ _15482_/X _15483_/X _15484_/X _24568_/Q _15466_/X VGND VGND VPWR VPWR _15485_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22436__B _22445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23676__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17224_ _11728_/C VGND VGND VPWR VPWR _17224_/Y sky130_fd_sc_hd__inv_2
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ _11647_/X VGND VGND VPWR VPWR _11648_/X sky130_fd_sc_hd__buf_2
X_14436_ _21403_/A _14436_/B VGND VGND VPWR VPWR _14437_/A sky130_fd_sc_hd__and2_4
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22155__C _22155_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17155_ _24032_/Q _17154_/Y VGND VGND VPWR VPWR _17156_/C sky130_fd_sc_hd__or2_4
X_11579_ _11579_/A VGND VGND VPWR VPWR _11579_/Y sky130_fd_sc_hd__inv_2
X_14367_ HREADY HSEL VGND VGND VPWR VPWR _14367_/Y sky130_fd_sc_hd__nand2_4
XFILLER_7_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14235__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16106_ _22232_/A _16099_/X _15978_/X _16105_/X VGND VGND VPWR VPWR _24333_/D sky130_fd_sc_hd__a2bb2o_4
X_13318_ _13222_/A _13314_/X _13318_/C VGND VGND VPWR VPWR _13318_/X sky130_fd_sc_hd__or3_4
XFILLER_115_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14298_ _14297_/Y _14293_/X _14221_/X _14293_/X VGND VGND VPWR VPWR _14298_/X sky130_fd_sc_hd__a2bb2o_4
X_17086_ _17086_/A VGND VGND VPWR VPWR _17086_/X sky130_fd_sc_hd__buf_2
XFILLER_6_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22452__A _20926_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16037_ _24355_/Q VGND VGND VPWR VPWR _16037_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13249_ _13146_/A _13249_/B VGND VGND VPWR VPWR _13249_/X sky130_fd_sc_hd__or2_4
XFILLER_131_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16450__A _16450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22171__B _22170_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16619__B1 _24125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21068__A _20926_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11594__A _16096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16634__A3 HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17988_ _22319_/A _17977_/X _15507_/X _17987_/X VGND VGND VPWR VPWR _23921_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24464__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19727_ _19709_/Y VGND VGND VPWR VPWR _19727_/X sky130_fd_sc_hd__buf_2
X_16939_ _16831_/D _16924_/B VGND VGND VPWR VPWR _16941_/B sky130_fd_sc_hd__nand2_4
XFILLER_38_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18377__A _18369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19658_ _23257_/Q VGND VGND VPWR VPWR _19658_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18609_ _23631_/Q _20279_/A VGND VGND VPWR VPWR _20283_/A sky130_fd_sc_hd__or2_4
X_19589_ _21383_/B _19588_/X _19459_/X _19588_/X VGND VGND VPWR VPWR _23281_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21620_ _17631_/Y _21611_/X _21619_/X VGND VGND VPWR VPWR _21620_/X sky130_fd_sc_hd__or3_4
XFILLER_52_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13314__A _13065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22340__A1 _24137_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19734__A2_N _19727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21551_ _14255_/Y _23025_/B _24788_/Q _21357_/X VGND VGND VPWR VPWR _21551_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20502_ _13509_/X _13497_/D VGND VGND VPWR VPWR _20502_/X sky130_fd_sc_hd__or2_4
X_24270_ _24104_/CLK _16272_/X HRESETn VGND VGND VPWR VPWR _22477_/A sky130_fd_sc_hd__dfrtp_4
X_21482_ _21935_/A _21482_/B VGND VGND VPWR VPWR _21482_/X sky130_fd_sc_hd__or2_4
XFILLER_105_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12872__B _21840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23221_ _23246_/CLK _23221_/D VGND VGND VPWR VPWR _23221_/Q sky130_fd_sc_hd__dfxtp_4
X_20433_ _13503_/X VGND VGND VPWR VPWR _20433_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23152_ _23135_/CLK _19942_/X VGND VGND VPWR VPWR _19941_/A sky130_fd_sc_hd__dfxtp_4
X_20364_ _20368_/B _20363_/Y _20349_/X VGND VGND VPWR VPWR _20364_/X sky130_fd_sc_hd__and3_4
XFILLER_49_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22103_ _20966_/A _22103_/B VGND VGND VPWR VPWR _22103_/X sky130_fd_sc_hd__or2_4
XFILLER_134_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15530__B1 _20413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23083_ _23109_/CLK _23083_/D VGND VGND VPWR VPWR _21795_/A sky130_fd_sc_hd__dfxtp_4
X_20295_ _20295_/A VGND VGND VPWR VPWR _23633_/D sky130_fd_sc_hd__inv_2
X_22034_ _20402_/A _21860_/B VGND VGND VPWR VPWR _22034_/X sky130_fd_sc_hd__and2_4
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19811__A3 _11643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17283__B1 _25200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14097__B1 _13645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24134__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21906__A1 _22806_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23985_ _23986_/CLK _17425_/X HRESETn VGND VGND VPWR VPWR _17257_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15704__A _11625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21425__B _21425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22936_ _13337_/A _22932_/Y _22407_/X _22935_/X VGND VGND VPWR VPWR _22936_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15597__B1 _24527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22867_ _22931_/A _22867_/B _22867_/C VGND VGND VPWR VPWR _22874_/C sky130_fd_sc_hd__and3_4
X_12620_ _25057_/Q VGND VGND VPWR VPWR _12701_/A sky130_fd_sc_hd__inv_2
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24606_ _24606_/CLK _15348_/X HRESETn VGND VGND VPWR VPWR _15347_/A sky130_fd_sc_hd__dfrtp_4
X_21818_ _20972_/A _19628_/Y VGND VGND VPWR VPWR _21818_/X sky130_fd_sc_hd__or2_4
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22798_ _15572_/A _22794_/X _20745_/X _22797_/X VGND VGND VPWR VPWR _22799_/A sky130_fd_sc_hd__o22a_4
XANTENNA__22537__A _21544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12551_ _12550_/X _24527_/Q _12549_/Y _24527_/Q VGND VGND VPWR VPWR _12552_/D sky130_fd_sc_hd__a2bb2o_4
X_21749_ _13428_/A _21400_/X _16393_/D _21748_/Y VGND VGND VPWR VPWR _21749_/X sky130_fd_sc_hd__a211o_4
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24537_ _23486_/CLK _24537_/D HRESETn VGND VGND VPWR VPWR _19828_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22882__A2 _21553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16535__A _16530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16010__A1 _15439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11502_ _11501_/X VGND VGND VPWR VPWR _11503_/A sky130_fd_sc_hd__buf_2
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12482_ _22564_/A _12481_/Y VGND VGND VPWR VPWR _12483_/C sky130_fd_sc_hd__or2_4
X_15270_ _15270_/A VGND VGND VPWR VPWR _15270_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24468_ _24488_/CLK _24468_/D HRESETn VGND VGND VPWR VPWR _12356_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14221_ _15282_/A VGND VGND VPWR VPWR _14221_/X sky130_fd_sc_hd__buf_2
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23419_ _23419_/CLK _23419_/D VGND VGND VPWR VPWR _23419_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14055__A _14055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24399_ _24399_/CLK _15901_/X HRESETn VGND VGND VPWR VPWR _15899_/A sky130_fd_sc_hd__dfrtp_4
X_14152_ _24838_/Q _14145_/X _14151_/Y VGND VGND VPWR VPWR _14152_/X sky130_fd_sc_hd__o21a_4
XFILLER_4_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13103_ _11741_/X VGND VGND VPWR VPWR _13182_/A sky130_fd_sc_hd__buf_2
X_14083_ _14083_/A VGND VGND VPWR VPWR _14083_/Y sky130_fd_sc_hd__inv_2
X_18960_ _18957_/Y _18958_/X _18959_/X _18958_/X VGND VGND VPWR VPWR _23505_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15521__B1 _24549_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24904__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13034_ _13050_/A _13032_/X _13033_/X VGND VGND VPWR VPWR _13034_/X sky130_fd_sc_hd__and3_4
X_17911_ _17879_/A _17909_/X _17911_/C VGND VGND VPWR VPWR _17911_/X sky130_fd_sc_hd__and3_4
X_18891_ _18876_/Y VGND VGND VPWR VPWR _18891_/X sky130_fd_sc_hd__buf_2
XFILLER_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17274__B1 _25195_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17842_ _17689_/X _17842_/B _17842_/C VGND VGND VPWR VPWR _17842_/X sky130_fd_sc_hd__and3_4
XANTENNA__21070__B2 _21069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17773_ _17879_/A _17770_/X _17772_/X VGND VGND VPWR VPWR _17777_/B sky130_fd_sc_hd__and3_4
XFILLER_134_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14985_ _14977_/C _14983_/X _14984_/X _14979_/B VGND VGND VPWR VPWR _14986_/A sky130_fd_sc_hd__a211o_4
X_19512_ _19508_/Y _19511_/X _19442_/X _19511_/X VGND VGND VPWR VPWR _19512_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16724_ _15970_/Y _22376_/A _15970_/Y _22376_/A VGND VGND VPWR VPWR _16726_/C sky130_fd_sc_hd__a2bb2o_4
X_13936_ _13936_/A VGND VGND VPWR VPWR _13937_/A sky130_fd_sc_hd__inv_2
XANTENNA__22570__A1 _22539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18774__B1 _18679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19443_ _19438_/Y _19441_/X _19442_/X _19441_/X VGND VGND VPWR VPWR _23334_/D sky130_fd_sc_hd__a2bb2o_4
X_16655_ _16655_/A VGND VGND VPWR VPWR _16655_/Y sky130_fd_sc_hd__inv_2
X_13867_ _13867_/A _13866_/Y _13867_/C _13830_/X VGND VGND VPWR VPWR _13868_/A sky130_fd_sc_hd__or4_4
XANTENNA__20581__B1 _20562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23857__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15606_ _12617_/Y _15604_/X _11563_/X _15604_/X VGND VGND VPWR VPWR _24522_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13134__A _13011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12818_ _25007_/Q VGND VGND VPWR VPWR _12818_/Y sky130_fd_sc_hd__inv_2
X_19374_ _19370_/Y _19373_/X _19329_/X _19373_/X VGND VGND VPWR VPWR _23358_/D sky130_fd_sc_hd__a2bb2o_4
X_16586_ _14833_/Y _16584_/X _16334_/X _16584_/X VGND VGND VPWR VPWR _16586_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13798_ _13798_/A VGND VGND VPWR VPWR _13798_/Y sky130_fd_sc_hd__inv_2
X_18325_ _18325_/A VGND VGND VPWR VPWR _18325_/Y sky130_fd_sc_hd__inv_2
X_15537_ _15558_/A VGND VGND VPWR VPWR _15537_/X sky130_fd_sc_hd__buf_2
X_12749_ _12749_/A _12742_/X _12749_/C VGND VGND VPWR VPWR _12749_/X sky130_fd_sc_hd__and3_4
XANTENNA__12973__A _21840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20884__A1 _12062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18256_ _18256_/A _18260_/B VGND VGND VPWR VPWR _18257_/C sky130_fd_sc_hd__or2_4
X_15468_ HWDATA[30] VGND VGND VPWR VPWR _15468_/X sky130_fd_sc_hd__buf_2
X_17207_ _17204_/Y _17198_/X _17205_/X _17206_/X VGND VGND VPWR VPWR _24017_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11589__A HWDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14419_ _14377_/B VGND VGND VPWR VPWR _14419_/Y sky130_fd_sc_hd__inv_2
X_18187_ _16048_/Y _23875_/Q _16048_/Y _23875_/Q VGND VGND VPWR VPWR _18190_/B sky130_fd_sc_hd__a2bb2o_4
X_15399_ _15398_/Y _15396_/X _15282_/X _15396_/X VGND VGND VPWR VPWR _24587_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17138_ _17028_/Y _17135_/X VGND VGND VPWR VPWR _17138_/X sky130_fd_sc_hd__or2_4
X_17069_ _24054_/Q _17074_/B VGND VGND VPWR VPWR _17069_/X sky130_fd_sc_hd__or2_4
XANTENNA__15512__B1 _15511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24645__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22389__B2 _20866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20080_ _21909_/B _20077_/X _19600_/A _20077_/X VGND VGND VPWR VPWR _20080_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19254__B2 _19251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13309__A _13309_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23770_ _24644_/CLK _20208_/Y HRESETn VGND VGND VPWR VPWR _23770_/Q sky130_fd_sc_hd__dfrtp_4
X_20982_ _22087_/A _20982_/B VGND VGND VPWR VPWR _20982_/X sky130_fd_sc_hd__or2_4
XANTENNA__18765__B1 _18764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22561__A1 _24412_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22721_ _21540_/X _22719_/X _20839_/X _22720_/X VGND VGND VPWR VPWR _22721_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20572__B1 _20562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22652_ _21064_/Y VGND VGND VPWR VPWR _22652_/X sky130_fd_sc_hd__buf_2
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14251__B1 _14232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22313__A1 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22313__B2 _22228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21603_ _17651_/A _19720_/Y VGND VGND VPWR VPWR _21603_/X sky130_fd_sc_hd__or2_4
XANTENNA__12262__C1 _12195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22583_ _16341_/A _22147_/X _22148_/X _22582_/X VGND VGND VPWR VPWR _22583_/X sky130_fd_sc_hd__a211o_4
XFILLER_55_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12883__A _12933_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21534_ _21534_/A _21402_/X VGND VGND VPWR VPWR _21534_/X sky130_fd_sc_hd__and2_4
X_24322_ _24071_/CLK _16130_/X HRESETn VGND VGND VPWR VPWR _16817_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24253_ _24222_/CLK _24253_/D HRESETn VGND VGND VPWR VPWR _16304_/A sky130_fd_sc_hd__dfrtp_4
X_21465_ _21461_/X _21464_/X _18049_/X VGND VGND VPWR VPWR _21465_/X sky130_fd_sc_hd__o21a_4
X_23204_ _24005_/CLK _19805_/X VGND VGND VPWR VPWR _23204_/Q sky130_fd_sc_hd__dfxtp_4
X_20416_ _20416_/A VGND VGND VPWR VPWR _20416_/X sky130_fd_sc_hd__buf_2
XFILLER_134_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24184_ _24185_/CLK _16491_/X HRESETn VGND VGND VPWR VPWR _24184_/Q sky130_fd_sc_hd__dfrtp_4
X_21396_ _21396_/A _21396_/B _21396_/C VGND VGND VPWR VPWR _21396_/X sky130_fd_sc_hd__or3_4
XFILLER_135_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23135_ _23135_/CLK _19987_/X VGND VGND VPWR VPWR _23135_/Q sky130_fd_sc_hd__dfxtp_4
X_20347_ _20347_/A VGND VGND VPWR VPWR _20347_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24386__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23066_ _24587_/CLK _20413_/A VGND VGND VPWR VPWR _23066_/Q sky130_fd_sc_hd__dfxtp_4
X_20278_ _18622_/X VGND VGND VPWR VPWR _20278_/X sky130_fd_sc_hd__buf_2
XFILLER_68_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15418__B _16475_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19245__B2 _19244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24315__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22017_ _22017_/A VGND VGND VPWR VPWR _22017_/X sky130_fd_sc_hd__buf_2
XFILLER_118_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_1_1_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11654__A2_N _23922_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_56_0_HCLK clkbuf_6_28_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_56_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11962__A _11961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14770_ _15044_/A VGND VGND VPWR VPWR _14770_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12096__A2 _24564_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11982_ _11980_/Y _11978_/X _11981_/X _11978_/X VGND VGND VPWR VPWR _25149_/D sky130_fd_sc_hd__a2bb2o_4
X_23968_ _23969_/CLK _23968_/D HRESETn VGND VGND VPWR VPWR _22853_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22552__B2 _22549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13721_ _13720_/X VGND VGND VPWR VPWR _13745_/D sky130_fd_sc_hd__inv_2
X_22919_ _22919_/A _22909_/X _22912_/X _22918_/X VGND VGND VPWR VPWR _22919_/X sky130_fd_sc_hd__or4_4
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23899_ _23898_/CLK _18056_/X HRESETn VGND VGND VPWR VPWR _21363_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23950__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16440_ _16438_/Y _16434_/X _15369_/X _16439_/X VGND VGND VPWR VPWR _16440_/X sky130_fd_sc_hd__a2bb2o_4
X_13652_ _13649_/A VGND VGND VPWR VPWR _13652_/X sky130_fd_sc_hd__buf_2
XANTENNA__25174__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14242__B1 _14221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22304__B2 _15824_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23801__D MSI_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12603_ _12730_/A VGND VGND VPWR VPWR _12731_/A sky130_fd_sc_hd__inv_2
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16371_ _16371_/A VGND VGND VPWR VPWR _16371_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25103__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13583_ _11673_/Y _13562_/X VGND VGND VPWR VPWR _13583_/Y sky130_fd_sc_hd__nand2_4
XFILLER_12_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15990__B1 _15897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18110_ _23885_/Q VGND VGND VPWR VPWR _18110_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15322_ _15322_/A _15531_/B VGND VGND VPWR VPWR _15325_/A sky130_fd_sc_hd__or2_4
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ _12534_/A _12537_/B VGND VGND VPWR VPWR _12534_/Y sky130_fd_sc_hd__nand2_4
X_19090_ _19088_/Y _19084_/X _19089_/X _19084_/X VGND VGND VPWR VPWR _23458_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18041_ _18022_/X _18061_/B _18039_/X VGND VGND VPWR VPWR _18041_/X sky130_fd_sc_hd__o21a_4
XFILLER_9_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15253_ _13769_/A _15247_/X _15240_/X _13761_/B _15245_/X VGND VGND VPWR VPWR _15253_/X
+ sky130_fd_sc_hd__a32o_4
X_12465_ _12489_/A _12465_/B _12464_/X VGND VGND VPWR VPWR _12466_/B sky130_fd_sc_hd__or3_4
XFILLER_138_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14204_ _24822_/Q VGND VGND VPWR VPWR _14204_/Y sky130_fd_sc_hd__inv_2
X_12396_ _12390_/X _12396_/B _12396_/C _12395_/X VGND VGND VPWR VPWR _12396_/X sky130_fd_sc_hd__or4_4
X_15184_ _14941_/Y _15159_/X _15126_/X _15182_/B VGND VGND VPWR VPWR _15184_/X sky130_fd_sc_hd__a211o_4
XANTENNA__20515__A _20465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14135_ _24845_/Q _14122_/X _24844_/Q _14127_/X VGND VGND VPWR VPWR _14135_/X sky130_fd_sc_hd__o22a_4
X_19992_ _19988_/Y _19991_/X _17993_/X _19991_/X VGND VGND VPWR VPWR _19992_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14066_ _13742_/D VGND VGND VPWR VPWR _14066_/Y sky130_fd_sc_hd__inv_2
X_18943_ _16035_/B _14592_/B _19144_/A VGND VGND VPWR VPWR _18943_/X sky130_fd_sc_hd__and3_4
XANTENNA__24056__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13017_ _13042_/A _13017_/B VGND VGND VPWR VPWR _13017_/X sky130_fd_sc_hd__or2_4
X_18874_ _18873_/X VGND VGND VPWR VPWR _18874_/X sky130_fd_sc_hd__buf_2
XFILLER_66_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17825_ _17924_/A _18771_/A VGND VGND VPWR VPWR _17827_/B sky130_fd_sc_hd__or2_4
XFILLER_121_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12968__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17756_ _14577_/X VGND VGND VPWR VPWR _17928_/A sky130_fd_sc_hd__buf_2
X_14968_ _24678_/Q _14956_/Y _15197_/A _24259_/Q VGND VGND VPWR VPWR _14972_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14481__B1 _14480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22543__A1 _12947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16707_ _16698_/X _16707_/B _16703_/X _16707_/D VGND VGND VPWR VPWR _16707_/X sky130_fd_sc_hd__or4_4
X_13919_ _13815_/X _20179_/C _13896_/X _13830_/C _13886_/X VGND VGND VPWR VPWR _13919_/X
+ sky130_fd_sc_hd__a32o_4
X_17687_ _17683_/X _17686_/X _14564_/X VGND VGND VPWR VPWR _17687_/X sky130_fd_sc_hd__o21a_4
X_14899_ _24660_/Q _14897_/Y _14898_/Y _24281_/Q VGND VGND VPWR VPWR _14905_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23691__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19426_ _19423_/Y _19418_/X _19424_/X _19425_/X VGND VGND VPWR VPWR _23340_/D sky130_fd_sc_hd__a2bb2o_4
X_16638_ _14781_/Y _16632_/X HWDATA[22] _16632_/X VGND VGND VPWR VPWR _24115_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14233__B1 _14232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23620__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21081__A _21113_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19357_ _13175_/B VGND VGND VPWR VPWR _19357_/Y sky130_fd_sc_hd__inv_2
X_16569_ _16575_/A VGND VGND VPWR VPWR _16570_/A sky130_fd_sc_hd__buf_2
XFILLER_52_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18308_ _18212_/Y _18311_/B _18228_/X VGND VGND VPWR VPWR _18308_/Y sky130_fd_sc_hd__a21oi_4
X_19288_ _19288_/A VGND VGND VPWR VPWR _21827_/B sky130_fd_sc_hd__inv_2
XFILLER_31_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24897__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18239_ _18239_/A VGND VGND VPWR VPWR _23873_/D sky130_fd_sc_hd__inv_2
XFILLER_102_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24826__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22624__B _22587_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21250_ _15428_/X VGND VGND VPWR VPWR _21250_/X sky130_fd_sc_hd__buf_2
XFILLER_135_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20425__A _20425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20201_ _20201_/A _20201_/B _20201_/C VGND VGND VPWR VPWR _20212_/D sky130_fd_sc_hd__or3_4
XANTENNA__16289__A1 _15915_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21181_ _21181_/A _21638_/A VGND VGND VPWR VPWR _21181_/X sky130_fd_sc_hd__or2_4
XANTENNA__21282__B2 _21562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20132_ _23077_/Q _20131_/Y _20709_/A _20131_/A VGND VGND VPWR VPWR _20132_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15500__A3 _15499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22607__A1_N _12412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20063_ _20062_/Y _20060_/X _15520_/X _20060_/X VGND VGND VPWR VPWR _23106_/D sky130_fd_sc_hd__a2bb2o_4
X_24940_ _24937_/CLK _24940_/D HRESETn VGND VGND VPWR VPWR _24940_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21585__A2 _22840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21256__A _20782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24871_ _24870_/CLK _14049_/X HRESETn VGND VGND VPWR VPWR _14045_/A sky130_fd_sc_hd__dfstp_4
XFILLER_85_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23779__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23822_ _23826_/CLK _23822_/D HRESETn VGND VGND VPWR VPWR _23822_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23708__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20965_ _20965_/A VGND VGND VPWR VPWR _20966_/A sky130_fd_sc_hd__buf_2
X_23753_ _23753_/CLK _20668_/X HRESETn VGND VGND VPWR VPWR _23753_/Q sky130_fd_sc_hd__dfrtp_4
X_22704_ _22364_/X _22703_/X _22634_/X _24523_/Q _22366_/X VGND VGND VPWR VPWR _22704_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_81_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21703__B _21703_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20896_ _20852_/Y _20868_/X _20878_/Y _20896_/D VGND VGND VPWR VPWR _20897_/A sky130_fd_sc_hd__or4_4
X_23684_ _24902_/CLK _23684_/D HRESETn VGND VGND VPWR VPWR _23684_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22635_ _22364_/X _22633_/X _22634_/X _24521_/Q _22366_/X VGND VGND VPWR VPWR _22635_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_110_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14775__B2 _14709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19163__B1 _19095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20848__B2 _21093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22566_ _24562_/Q _22557_/X _20800_/X _22565_/X VGND VGND VPWR VPWR _22566_/X sky130_fd_sc_hd__a211o_4
XFILLER_22_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21517_ _21385_/A _21517_/B VGND VGND VPWR VPWR _21519_/B sky130_fd_sc_hd__or2_4
X_24305_ _24037_/CLK _24305_/D HRESETn VGND VGND VPWR VPWR _24305_/Q sky130_fd_sc_hd__dfrtp_4
X_22497_ _16515_/Y _22497_/B VGND VGND VPWR VPWR _22497_/X sky130_fd_sc_hd__and2_4
XFILLER_33_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16813__A _17053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24567__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12250_ _12237_/X VGND VGND VPWR VPWR _12250_/Y sky130_fd_sc_hd__inv_2
X_21448_ _24917_/Q _21448_/B VGND VGND VPWR VPWR _21448_/X sky130_fd_sc_hd__and2_4
X_24236_ _24201_/CLK _24236_/D HRESETn VGND VGND VPWR VPWR _24236_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11957__A _15422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12181_ _12176_/X _12178_/X _12180_/X VGND VGND VPWR VPWR _12256_/B sky130_fd_sc_hd__or3_4
XANTENNA__22470__B1 _24560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24167_ _24167_/CLK _16533_/X HRESETn VGND VGND VPWR VPWR _16532_/A sky130_fd_sc_hd__dfrtp_4
X_21379_ _21394_/A _21377_/X _21379_/C VGND VGND VPWR VPWR _21379_/X sky130_fd_sc_hd__and3_4
XFILLER_123_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23068__D HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23118_ _23293_/CLK _20032_/X VGND VGND VPWR VPWR _23118_/Q sky130_fd_sc_hd__dfxtp_4
X_24098_ _24098_/CLK _24098_/D HRESETn VGND VGND VPWR VPWR _24098_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21025__A1 _20940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15940_ _22783_/A VGND VGND VPWR VPWR _15940_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23049_ VGND VGND VPWR VPWR _23049_/HI scl_o_S5 sky130_fd_sc_hd__conb_1
XFILLER_27_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15871_ _15870_/Y _15868_/X _11581_/X _15868_/X VGND VGND VPWR VPWR _15871_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17610_ _17603_/A _17594_/B _17609_/X VGND VGND VPWR VPWR _23947_/D sky130_fd_sc_hd__and3_4
X_14822_ _24691_/Q _14821_/A _14743_/X _14821_/Y VGND VGND VPWR VPWR _14822_/X sky130_fd_sc_hd__o22a_4
XFILLER_95_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18590_ _16368_/Y _23820_/Q _16368_/Y _23820_/Q VGND VGND VPWR VPWR _18590_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18729__B1 _18685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17541_ _17532_/X VGND VGND VPWR VPWR _17545_/B sky130_fd_sc_hd__inv_2
X_14753_ _24699_/Q _14751_/Y _14869_/B _24098_/Q VGND VGND VPWR VPWR _14753_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11965_ _22982_/A _11956_/X VGND VGND VPWR VPWR _11965_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__20536__B1 _20511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13704_ _24916_/Q _13686_/X _24915_/Q _13681_/X VGND VGND VPWR VPWR _13704_/X sky130_fd_sc_hd__o22a_4
XFILLER_45_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_143_0_HCLK clkbuf_7_71_0_HCLK/X VGND VGND VPWR VPWR _25061_/CLK sky130_fd_sc_hd__clkbuf_1
X_17472_ _21801_/A _17457_/B VGND VGND VPWR VPWR _17472_/X sky130_fd_sc_hd__or2_4
X_14684_ _14680_/Y _14683_/Y _14676_/X VGND VGND VPWR VPWR _14684_/X sky130_fd_sc_hd__o21a_4
X_11896_ _20688_/A VGND VGND VPWR VPWR _11896_/Y sky130_fd_sc_hd__inv_2
X_19211_ _22046_/A VGND VGND VPWR VPWR _19211_/Y sky130_fd_sc_hd__inv_2
X_16423_ _24210_/Q VGND VGND VPWR VPWR _16423_/Y sky130_fd_sc_hd__inv_2
X_13635_ _15282_/A VGND VGND VPWR VPWR _13635_/X sky130_fd_sc_hd__buf_2
XANTENNA__22289__B1 _14709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19154__B1 _19152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19142_ _19141_/Y _19137_/X _19120_/X _19137_/A VGND VGND VPWR VPWR _23439_/D sky130_fd_sc_hd__a2bb2o_4
X_16354_ _16354_/A VGND VGND VPWR VPWR _16354_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13566_ _11653_/A _13566_/B _13566_/C _13566_/D VGND VGND VPWR VPWR _13567_/A sky130_fd_sc_hd__and4_4
XANTENNA__24990__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15305_ _15314_/B _15301_/X HADDR[22] _15304_/X VGND VGND VPWR VPWR _15305_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14518__A1 _14506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12517_ _12345_/X _12515_/X _12516_/Y VGND VGND VPWR VPWR _25079_/D sky130_fd_sc_hd__o21a_4
X_19073_ _23464_/Q VGND VGND VPWR VPWR _19073_/Y sky130_fd_sc_hd__inv_2
X_16285_ _14887_/Y _16282_/X _15894_/X _16282_/X VGND VGND VPWR VPWR _16285_/X sky130_fd_sc_hd__a2bb2o_4
X_13497_ _20512_/A _20513_/B _23717_/Q _13497_/D VGND VGND VPWR VPWR _13510_/B sky130_fd_sc_hd__or4_4
XFILLER_121_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22444__B _22444_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18024_ _18023_/X VGND VGND VPWR VPWR _18025_/D sky130_fd_sc_hd__buf_2
X_15236_ _15236_/A _15235_/Y VGND VGND VPWR VPWR _15237_/B sky130_fd_sc_hd__or2_4
X_12448_ _12448_/A _12448_/B VGND VGND VPWR VPWR _12451_/B sky130_fd_sc_hd__or2_4
XFILLER_138_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24237__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21264__A1 _22501_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_5_11_0_HCLK_A clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15167_ _15166_/X VGND VGND VPWR VPWR _24670_/D sky130_fd_sc_hd__inv_2
XFILLER_114_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12379_ _21566_/A VGND VGND VPWR VPWR _12379_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14118_ _14107_/Y _14116_/X _14117_/Y VGND VGND VPWR VPWR _14118_/X sky130_fd_sc_hd__o21a_4
X_15098_ _15158_/A VGND VGND VPWR VPWR _15154_/A sky130_fd_sc_hd__buf_2
X_19975_ _19982_/A VGND VGND VPWR VPWR _19975_/X sky130_fd_sc_hd__buf_2
XANTENNA__17554__A _16692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22213__B1 _21886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14049_ _14045_/Y _14048_/X _13663_/X _14048_/X VGND VGND VPWR VPWR _14049_/X sky130_fd_sc_hd__a2bb2o_4
X_18926_ _18926_/A VGND VGND VPWR VPWR _18926_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16691__B2 _22853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22764__A1 _21572_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18857_ _18856_/Y _18854_/X _18740_/X _18854_/X VGND VGND VPWR VPWR _18857_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15246__A2 _14100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23872__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17808_ _17878_/A _17808_/B VGND VGND VPWR VPWR _17809_/C sky130_fd_sc_hd__or2_4
X_18788_ _18787_/Y _18785_/X _18740_/X _18785_/X VGND VGND VPWR VPWR _23565_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25096__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21319__A2 _11514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22516__A1 _22116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22516__B2 _22118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23801__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17739_ _17739_/A _17739_/B _17739_/C VGND VGND VPWR VPWR _17739_/X sky130_fd_sc_hd__and3_4
XANTENNA__25025__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19393__B1 _19392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20750_ _20749_/X VGND VGND VPWR VPWR _20750_/X sky130_fd_sc_hd__buf_2
XFILLER_35_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19409_ _19396_/Y VGND VGND VPWR VPWR _19409_/X sky130_fd_sc_hd__buf_2
X_20681_ _20679_/Y _20680_/Y _13543_/B VGND VGND VPWR VPWR _20681_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15954__B1 _15772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22420_ _22420_/A _22147_/A VGND VGND VPWR VPWR _22420_/X sky130_fd_sc_hd__and2_4
XFILLER_17_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22351_ _22351_/A VGND VGND VPWR VPWR _22351_/X sky130_fd_sc_hd__buf_2
XANTENNA__24660__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21302_ _21570_/A _21302_/B _21302_/C VGND VGND VPWR VPWR _21323_/A sky130_fd_sc_hd__and3_4
X_25070_ _25091_/CLK _12539_/X HRESETn VGND VGND VPWR VPWR _12322_/A sky130_fd_sc_hd__dfrtp_4
X_22282_ _22282_/A _22281_/X VGND VGND VPWR VPWR _22282_/X sky130_fd_sc_hd__and2_4
XANTENNA__20871__A2_N _21638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24021_ _23668_/CLK _24021_/D HRESETn VGND VGND VPWR VPWR _20723_/B sky130_fd_sc_hd__dfstp_4
X_21233_ _21227_/A _21233_/B VGND VGND VPWR VPWR _21233_/X sky130_fd_sc_hd__or2_4
XFILLER_85_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21164_ _21348_/A _19703_/Y VGND VGND VPWR VPWR _21167_/B sky130_fd_sc_hd__or2_4
XFILLER_104_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20115_ _20982_/B _20110_/X _25169_/Q _20110_/A VGND VGND VPWR VPWR _23086_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21095_ _22017_/A _21094_/X VGND VGND VPWR VPWR _21095_/X sky130_fd_sc_hd__or2_4
XFILLER_63_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21558__A2 _21553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20046_ _21475_/B _20041_/X _19724_/X _20041_/X VGND VGND VPWR VPWR _20046_/X sky130_fd_sc_hd__a2bb2o_4
X_24923_ _24923_/CLK _24923_/D HRESETn VGND VGND VPWR VPWR _20201_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19620__B2 _19613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24854_ _24728_/CLK _24854_/D HRESETn VGND VGND VPWR VPWR _23655_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_27_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23805_ _24897_/CLK _23805_/D HRESETn VGND VGND VPWR VPWR _20715_/A sky130_fd_sc_hd__dfrtp_4
X_24785_ _24776_/CLK _24785_/D HRESETn VGND VGND VPWR VPWR _24785_/Q sky130_fd_sc_hd__dfrtp_4
X_21997_ _20747_/X _21989_/Y _21991_/X _21996_/X VGND VGND VPWR VPWR _21997_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11749_/X _11733_/B _11737_/Y VGND VGND VPWR VPWR _11761_/B sky130_fd_sc_hd__o21a_4
XPHY_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23736_ _24167_/CLK _20597_/Y HRESETn VGND VGND VPWR VPWR _23736_/Q sky130_fd_sc_hd__dfrtp_4
X_20948_ _22089_/A _20945_/X _20947_/X VGND VGND VPWR VPWR _20948_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_216_0_HCLK clkbuf_7_108_0_HCLK/X VGND VGND VPWR VPWR _24244_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11679_/A _23918_/Q _11679_/Y _11680_/Y VGND VGND VPWR VPWR _11681_/X sky130_fd_sc_hd__o22a_4
XFILLER_14_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23667_ _24723_/CLK _20347_/Y HRESETn VGND VGND VPWR VPWR _20345_/A sky130_fd_sc_hd__dfrtp_4
X_20879_ _22859_/A VGND VGND VPWR VPWR _22311_/A sky130_fd_sc_hd__buf_2
XANTENNA__21740__A1_N _14234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24748__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13419_/Y _14420_/A _13419_/Y _14420_/A VGND VGND VPWR VPWR _13420_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22618_ _24144_/Q _15692_/A _22576_/X _22617_/X VGND VGND VPWR VPWR _22619_/C sky130_fd_sc_hd__a211o_4
XPHY_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23598_ _25009_/CLK _23598_/D VGND VGND VPWR VPWR _23598_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13351_ _13338_/Y VGND VGND VPWR VPWR _13351_/X sky130_fd_sc_hd__buf_2
XANTENNA__21494__B2 _12063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24810__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22549_ _22549_/A VGND VGND VPWR VPWR _22549_/X sky130_fd_sc_hd__buf_2
XFILLER_122_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12302_ _12302_/A VGND VGND VPWR VPWR _12302_/Y sky130_fd_sc_hd__inv_2
X_16070_ _24345_/Q VGND VGND VPWR VPWR _16070_/Y sky130_fd_sc_hd__inv_2
X_13282_ _13065_/X _13280_/X _13281_/X VGND VGND VPWR VPWR _13282_/X sky130_fd_sc_hd__and3_4
XANTENNA__16370__B1 _16369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24330__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15021_ _14877_/D _15020_/X VGND VGND VPWR VPWR _15021_/X sky130_fd_sc_hd__or2_4
X_12233_ _12175_/A _12230_/X VGND VGND VPWR VPWR _12233_/X sky130_fd_sc_hd__or2_4
XANTENNA__15159__A _15159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24219_ _24192_/CLK _24219_/D HRESETn VGND VGND VPWR VPWR _24219_/Q sky130_fd_sc_hd__dfrtp_4
X_25199_ _23957_/CLK _11605_/X HRESETn VGND VGND VPWR VPWR _25199_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22994__A1 _21864_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12164_ _12423_/A VGND VGND VPWR VPWR _12418_/C sky130_fd_sc_hd__buf_2
XANTENNA__16122__B1 _15801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22280__A _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12095_ _24564_/Q VGND VGND VPWR VPWR _12095_/Y sky130_fd_sc_hd__inv_2
X_16972_ _16965_/X _16972_/B _16972_/C _16972_/D VGND VGND VPWR VPWR _16972_/X sky130_fd_sc_hd__or4_4
X_19760_ _19759_/Y VGND VGND VPWR VPWR _19760_/X sky130_fd_sc_hd__buf_2
XFILLER_96_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22746__A1 _24278_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15923_ _15922_/X VGND VGND VPWR VPWR _15923_/X sky130_fd_sc_hd__buf_2
X_18711_ _13644_/A VGND VGND VPWR VPWR _18711_/X sky130_fd_sc_hd__buf_2
XFILLER_42_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19691_ _23245_/Q VGND VGND VPWR VPWR _19691_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18642_ _14544_/A _14452_/X _14482_/X VGND VGND VPWR VPWR _19883_/C sky130_fd_sc_hd__or3_4
X_15854_ _15847_/A VGND VGND VPWR VPWR _15854_/X sky130_fd_sc_hd__buf_2
XFILLER_91_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_26_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_26_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14805_ _14798_/X _14799_/X _14802_/X _14804_/X VGND VGND VPWR VPWR _14805_/X sky130_fd_sc_hd__or4_4
XFILLER_64_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18573_ _16312_/A _23842_/Q _16312_/Y _18412_/A VGND VGND VPWR VPWR _18573_/X sky130_fd_sc_hd__o22a_4
X_15785_ _15781_/X _15582_/A _15505_/X _22365_/A _15779_/X VGND VGND VPWR VPWR _24441_/D
+ sky130_fd_sc_hd__a32o_4
X_12997_ _12996_/X VGND VGND VPWR VPWR _12997_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16718__A _16718_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17524_ _17524_/A VGND VGND VPWR VPWR _17524_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22439__B _22439_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14736_ _14876_/C VGND VGND VPWR VPWR _14736_/X sky130_fd_sc_hd__buf_2
X_11948_ _24620_/Q VGND VGND VPWR VPWR _11949_/A sky130_fd_sc_hd__buf_2
XANTENNA__16189__B1 _16096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17455_ _21799_/A VGND VGND VPWR VPWR _17455_/Y sky130_fd_sc_hd__inv_2
X_14667_ _24721_/Q _14610_/X _24721_/Q _14610_/X VGND VGND VPWR VPWR _14667_/X sky130_fd_sc_hd__a2bb2o_4
X_11879_ _11879_/A VGND VGND VPWR VPWR _22030_/A sky130_fd_sc_hd__inv_2
XANTENNA__24489__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16406_ _24217_/Q VGND VGND VPWR VPWR _16406_/Y sky130_fd_sc_hd__inv_2
X_13618_ _13618_/A VGND VGND VPWR VPWR _16305_/A sky130_fd_sc_hd__buf_2
XANTENNA__12859__A2_N _24432_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17386_ _17270_/Y _17386_/B VGND VGND VPWR VPWR _17386_/X sky130_fd_sc_hd__or2_4
X_14598_ _14597_/X VGND VGND VPWR VPWR _14598_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24418__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19125_ _19137_/A VGND VGND VPWR VPWR _19125_/X sky130_fd_sc_hd__buf_2
X_16337_ _16336_/Y _16333_/X _16259_/X _16333_/X VGND VGND VPWR VPWR _16337_/X sky130_fd_sc_hd__a2bb2o_4
X_13549_ _13549_/A VGND VGND VPWR VPWR _13549_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19056_ _14581_/Y _19123_/B VGND VGND VPWR VPWR _19100_/B sky130_fd_sc_hd__or2_4
X_16268_ _16228_/A VGND VGND VPWR VPWR _16268_/X sky130_fd_sc_hd__buf_2
XANTENNA__24071__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18007_ _18007_/A VGND VGND VPWR VPWR _18007_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20667__B1_N _13539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15219_ _15219_/A _15219_/B _15226_/C VGND VGND VPWR VPWR _24655_/D sky130_fd_sc_hd__and3_4
XANTENNA__11597__A HWDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16199_ _16198_/Y _16196_/X _15982_/X _16196_/X VGND VGND VPWR VPWR _24297_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24000__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22985__A1 _24155_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16113__B1 _15894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22190__A _22163_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20703__A scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15467__A2 _15461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19958_ _19957_/Y _19953_/X _15522_/X _19953_/X VGND VGND VPWR VPWR _23146_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_108_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_108_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22737__A1 _24567_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18909_ _18908_/Y _18906_/X _18817_/X _18906_/X VGND VGND VPWR VPWR _23523_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25206__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19889_ _23172_/Q VGND VGND VPWR VPWR _21784_/B sky130_fd_sc_hd__inv_2
XFILLER_83_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12150__B2 _24565_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21920_ _21342_/A _19762_/Y VGND VGND VPWR VPWR _21920_/X sky130_fd_sc_hd__or2_4
X_21851_ _21851_/A _20786_/A VGND VGND VPWR VPWR _21851_/X sky130_fd_sc_hd__or2_4
XFILLER_23_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20802_ _20759_/X VGND VGND VPWR VPWR _20802_/X sky130_fd_sc_hd__buf_2
XFILLER_58_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21782_ _21224_/A _21780_/X _21781_/X VGND VGND VPWR VPWR _21782_/X sky130_fd_sc_hd__and3_4
XFILLER_64_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24570_ _24488_/CLK _24570_/D HRESETn VGND VGND VPWR VPWR _24570_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21173__B1 _21172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23521_ _23560_/CLK _18914_/X VGND VGND VPWR VPWR _23521_/Q sky130_fd_sc_hd__dfxtp_4
X_20733_ _20733_/A _20733_/B VGND VGND VPWR VPWR _20733_/Y sky130_fd_sc_hd__nor2_4
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20920__B1 _20918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19118__B1 _19095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24841__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20664_ _23752_/Q _23751_/Q _20660_/B VGND VGND VPWR VPWR _20664_/X sky130_fd_sc_hd__or3_4
XFILLER_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23452_ _23440_/CLK _19107_/X VGND VGND VPWR VPWR _23452_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24159__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_46_0_HCLK clkbuf_8_47_0_HCLK/A VGND VGND VPWR VPWR _23560_/CLK sky130_fd_sc_hd__clkbuf_1
X_22403_ _22225_/X _22400_/X _22231_/X _22402_/X VGND VGND VPWR VPWR _22404_/B sky130_fd_sc_hd__o22a_4
XFILLER_137_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17459__A _21491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23383_ _23383_/CLK _19301_/X VGND VGND VPWR VPWR _19300_/A sky130_fd_sc_hd__dfxtp_4
X_20595_ _20594_/Y _20590_/Y _13534_/B VGND VGND VPWR VPWR _20595_/X sky130_fd_sc_hd__o21a_4
XFILLER_13_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12891__A _12921_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25122_ _24573_/CLK _12236_/Y HRESETn VGND VGND VPWR VPWR _25122_/Q sky130_fd_sc_hd__dfrtp_4
X_22334_ _22334_/A VGND VGND VPWR VPWR _22691_/A sky130_fd_sc_hd__buf_2
XFILLER_124_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22265_ _14897_/Y _22265_/B VGND VGND VPWR VPWR _22265_/X sky130_fd_sc_hd__and2_4
XFILLER_30_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25053_ _24521_/CLK _12720_/X HRESETn VGND VGND VPWR VPWR _25053_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22976__A1 _16621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21216_ _14524_/A _21214_/X _21215_/X VGND VGND VPWR VPWR _21216_/X sky130_fd_sc_hd__and3_4
XANTENNA__22976__B2 _21694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24004_ _25217_/CLK _24004_/D HRESETn VGND VGND VPWR VPWR _24004_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21709__A _21434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22196_ _16195_/A _20757_/A VGND VGND VPWR VPWR _22196_/X sky130_fd_sc_hd__or2_4
XFILLER_105_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23794__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21147_ _21147_/A _21145_/X _21146_/X VGND VGND VPWR VPWR _21147_/X sky130_fd_sc_hd__and3_4
XFILLER_133_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22728__B2 _22549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23723__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14130__A2 _14122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21078_ _21077_/X VGND VGND VPWR VPWR _21078_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12920_ _12781_/Y _12920_/B VGND VGND VPWR VPWR _12920_/X sky130_fd_sc_hd__or2_4
X_20029_ _20029_/A VGND VGND VPWR VPWR _21134_/B sky130_fd_sc_hd__inv_2
XFILLER_115_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17922__A _17725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24906_ _24904_/CLK _24906_/D HRESETn VGND VGND VPWR VPWR _24906_/Q sky130_fd_sc_hd__dfrtp_4
X_12851_ _24449_/Q VGND VGND VPWR VPWR _12851_/Y sky130_fd_sc_hd__inv_2
X_24837_ _24840_/CLK _24837_/D HRESETn VGND VGND VPWR VPWR _18111_/B sky130_fd_sc_hd__dfstp_4
XFILLER_41_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17245__A2_N _17415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24929__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11802_ _11802_/A _11801_/X _11802_/C VGND VGND VPWR VPWR _11803_/B sky130_fd_sc_hd__and3_4
X_15570_ _21292_/A VGND VGND VPWR VPWR _22884_/B sky130_fd_sc_hd__buf_2
X_12782_ _12781_/Y _24454_/Q _12781_/Y _24454_/Q VGND VGND VPWR VPWR _12782_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24768_ _24968_/CLK _14389_/X HRESETn VGND VGND VPWR VPWR _24768_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14521_ _21534_/A _14437_/X _14476_/Y VGND VGND VPWR VPWR _14521_/X sky130_fd_sc_hd__o21a_4
XPHY_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11733_ _11733_/A _11733_/B VGND VGND VPWR VPWR _11733_/X sky130_fd_sc_hd__and2_4
XPHY_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23719_ _23753_/CLK _20526_/X HRESETn VGND VGND VPWR VPWR _20524_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24582__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24699_ _24706_/CLK _24699_/D HRESETn VGND VGND VPWR VPWR _24699_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17240_ _11614_/A _17317_/D _11539_/Y _17352_/A VGND VGND VPWR VPWR _17242_/C sky130_fd_sc_hd__a2bb2o_4
XPHY_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _24739_/Q VGND VGND VPWR VPWR _14452_/X sky130_fd_sc_hd__buf_2
XFILLER_109_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11663_/Y _23913_/Q _11663_/Y _23913_/Q VGND VGND VPWR VPWR _11664_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22275__A _21581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24511__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _13403_/A VGND VGND VPWR VPWR _13403_/Y sky130_fd_sc_hd__inv_2
XPHY_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17171_ _17170_/Y VGND VGND VPWR VPWR _17171_/X sky130_fd_sc_hd__buf_2
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14383_ _14383_/A _14383_/B VGND VGND VPWR VPWR _14402_/B sky130_fd_sc_hd__or2_4
X_11595_ _11592_/Y _11588_/X _11594_/X _11588_/X VGND VGND VPWR VPWR _11595_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16122_ _16121_/Y _16117_/X _15801_/X _16117_/X VGND VGND VPWR VPWR _16122_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13334_ _20818_/A VGND VGND VPWR VPWR _13334_/X sky130_fd_sc_hd__buf_2
XFILLER_128_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16053_ _16050_/Y _16046_/X _15753_/X _16052_/X VGND VGND VPWR VPWR _16053_/X sky130_fd_sc_hd__a2bb2o_4
X_13265_ _13297_/A _23070_/Q VGND VGND VPWR VPWR _13267_/B sky130_fd_sc_hd__or2_4
X_15004_ _15004_/A _15012_/A VGND VGND VPWR VPWR _15014_/B sky130_fd_sc_hd__or2_4
XANTENNA__22967__A1 _15463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12904__B1 _12896_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12216_ _12219_/A _12219_/B VGND VGND VPWR VPWR _12216_/X sky130_fd_sc_hd__or2_4
XANTENNA__22967__B2 _22576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13196_ _13122_/A _13194_/X _13195_/X VGND VGND VPWR VPWR _13196_/X sky130_fd_sc_hd__and3_4
X_19812_ _19812_/A VGND VGND VPWR VPWR _22072_/B sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0_HCLK_A HCLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12147_ _12185_/B _24571_/Q _25122_/Q _12146_/Y VGND VGND VPWR VPWR _12147_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22719__B2 _22537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19743_ _19737_/Y VGND VGND VPWR VPWR _19743_/X sky130_fd_sc_hd__buf_2
X_12078_ _12078_/A VGND VGND VPWR VPWR _12078_/Y sky130_fd_sc_hd__inv_2
X_16955_ _24060_/Q _16954_/Y VGND VGND VPWR VPWR _16955_/X sky130_fd_sc_hd__or2_4
XFILLER_42_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12153__A2_N _24548_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15906_ _24396_/Q VGND VGND VPWR VPWR _15906_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17832__A _17725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16886_ _16800_/Y _16885_/X VGND VGND VPWR VPWR _16887_/A sky130_fd_sc_hd__or2_4
X_19674_ _19672_/Y _19668_/X _19603_/X _19673_/X VGND VGND VPWR VPWR _19674_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15837_ HWDATA[28] VGND VGND VPWR VPWR _15837_/X sky130_fd_sc_hd__buf_2
X_18625_ _18607_/X _18621_/X _23810_/Q _23811_/Q _18624_/X VGND VGND VPWR VPWR _18625_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_18_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21073__B _21113_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15768_ _15767_/X VGND VGND VPWR VPWR _15768_/X sky130_fd_sc_hd__buf_2
X_18556_ _18484_/A _18552_/X _18555_/Y VGND VGND VPWR VPWR _23815_/D sky130_fd_sc_hd__and3_4
XFILLER_79_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14719_ _14708_/X _14719_/B _14719_/C _14718_/X VGND VGND VPWR VPWR _14750_/B sky130_fd_sc_hd__or4_4
X_17507_ _23012_/A _17508_/B VGND VGND VPWR VPWR _17509_/B sky130_fd_sc_hd__or2_4
X_18487_ _18434_/X _18495_/D VGND VGND VPWR VPWR _18488_/B sky130_fd_sc_hd__or2_4
XANTENNA__15909__B1 _15291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15699_ _12329_/Y _15695_/X _15513_/X _15698_/X VGND VGND VPWR VPWR _15699_/X sky130_fd_sc_hd__a2bb2o_4
X_17438_ _17438_/A _17438_/B _17428_/C VGND VGND VPWR VPWR _17438_/X sky130_fd_sc_hd__and3_4
XANTENNA__16582__B1 _24148_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24252__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_5_0_HCLK clkbuf_8_5_0_HCLK/A VGND VGND VPWR VPWR _25183_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_119_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17369_ _17368_/X VGND VGND VPWR VPWR _24000_/D sky130_fd_sc_hd__inv_2
XFILLER_119_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20417__B _13517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19108_ _17807_/B VGND VGND VPWR VPWR _19108_/Y sky130_fd_sc_hd__inv_2
X_20380_ _20380_/A VGND VGND VPWR VPWR _20380_/Y sky130_fd_sc_hd__inv_2
X_19039_ _19037_/Y _19035_/X _19038_/X _19035_/X VGND VGND VPWR VPWR _23477_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22958__A1 _24574_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22050_ _22045_/X _22049_/X _20820_/X VGND VGND VPWR VPWR _22050_/X sky130_fd_sc_hd__o21a_4
XFILLER_86_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21529__A _21245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20969__B1 _20968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21001_ _20998_/A _21001_/B VGND VGND VPWR VPWR _21001_/X sky130_fd_sc_hd__or2_4
XFILLER_88_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16637__B2 _16622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15527__A _15418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25040__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12123__B2 _24550_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17742__A _17742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22952_ _24056_/Q _22952_/B VGND VGND VPWR VPWR _22955_/B sky130_fd_sc_hd__or2_4
XFILLER_112_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21903_ _17201_/Y _22153_/B _23660_/Q _21088_/X VGND VGND VPWR VPWR _21905_/C sky130_fd_sc_hd__a2bb2o_4
X_22883_ _22883_/A _20807_/X VGND VGND VPWR VPWR _22883_/X sky130_fd_sc_hd__and2_4
XFILLER_83_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19339__B1 _19201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24622_ _24587_/CLK _15303_/X HRESETn VGND VGND VPWR VPWR _24622_/Q sky130_fd_sc_hd__dfrtp_4
X_21834_ _22089_/A _21830_/X _21831_/X _21832_/X _21833_/X VGND VGND VPWR VPWR _21834_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_55_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24553_ _24566_/CLK _15515_/X HRESETn VGND VGND VPWR VPWR _12098_/A sky130_fd_sc_hd__dfrtp_4
X_21765_ _21760_/X _19447_/Y VGND VGND VPWR VPWR _21767_/B sky130_fd_sc_hd__or2_4
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23504_ _23511_/CLK _23504_/D VGND VGND VPWR VPWR _17935_/B sky130_fd_sc_hd__dfxtp_4
X_20716_ sda_oen_o_S4 _24769_/Q _20710_/A _13864_/X _20715_/Y VGND VGND VPWR VPWR
+ _20716_/X sky130_fd_sc_hd__a32o_4
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24484_ _24488_/CLK _15683_/X HRESETn VGND VGND VPWR VPWR _22565_/A sky130_fd_sc_hd__dfrtp_4
X_21696_ _21696_/A _21251_/A VGND VGND VPWR VPWR _21696_/X sky130_fd_sc_hd__and2_4
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23435_ _25067_/CLK _23435_/D VGND VGND VPWR VPWR _19155_/A sky130_fd_sc_hd__dfxtp_4
X_20647_ _20647_/A VGND VGND VPWR VPWR _20647_/X sky130_fd_sc_hd__buf_2
XFILLER_71_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16093__A _16093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14606__A _23665_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20578_ _20578_/A VGND VGND VPWR VPWR _20578_/Y sky130_fd_sc_hd__inv_2
X_23366_ _23374_/CLK _19351_/X VGND VGND VPWR VPWR _13017_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23975__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25105_ _25112_/CLK _12295_/X HRESETn VGND VGND VPWR VPWR _12152_/A sky130_fd_sc_hd__dfrtp_4
X_22317_ _22263_/X _22317_/B VGND VGND VPWR VPWR _22317_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__25199__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23297_ _23401_/CLK _19547_/X VGND VGND VPWR VPWR _19545_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22949__B2 _22549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23904__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13050_ _13050_/A _13048_/X _13050_/C VGND VGND VPWR VPWR _13050_/X sky130_fd_sc_hd__and3_4
X_25036_ _24435_/CLK _25036_/D HRESETn VGND VGND VPWR VPWR _23013_/A sky130_fd_sc_hd__dfrtp_4
X_22248_ _22248_/A VGND VGND VPWR VPWR _22248_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25128__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12001_ _12001_/A VGND VGND VPWR VPWR _12001_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11965__A _22982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22179_ _12098_/Y _21178_/A _12329_/Y _22228_/A VGND VGND VPWR VPWR _22180_/B sky130_fd_sc_hd__o22a_4
XFILLER_121_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16740_ _15995_/Y _23945_/Q _21044_/A _17614_/A VGND VGND VPWR VPWR _16740_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13952_ _13952_/A VGND VGND VPWR VPWR _13952_/X sky130_fd_sc_hd__buf_2
XFILLER_101_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12903_ _12921_/A _12901_/X _12902_/X VGND VGND VPWR VPWR _25034_/D sky130_fd_sc_hd__and3_4
XANTENNA__21174__A _17636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16671_ _16291_/A VGND VGND VPWR VPWR _16671_/X sky130_fd_sc_hd__buf_2
X_13883_ _13885_/A VGND VGND VPWR VPWR _13905_/A sky130_fd_sc_hd__buf_2
XFILLER_62_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16268__A _16228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24763__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15622_ _12556_/Y _15621_/X _13658_/X _15621_/X VGND VGND VPWR VPWR _24512_/D sky130_fd_sc_hd__a2bb2o_4
X_18410_ _18484_/A VGND VGND VPWR VPWR _18463_/A sky130_fd_sc_hd__buf_2
X_12834_ _12833_/X _22420_/A _12833_/X _22420_/A VGND VGND VPWR VPWR _12835_/D sky130_fd_sc_hd__a2bb2o_4
X_19390_ _19389_/Y _19386_/X _19366_/X _19386_/X VGND VGND VPWR VPWR _23352_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21324__D _21323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18341_ _16389_/Y _18442_/A _16389_/Y _23844_/Q VGND VGND VPWR VPWR _18347_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18002__B1 _16671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15553_ _19455_/A VGND VGND VPWR VPWR _15553_/Y sky130_fd_sc_hd__inv_2
X_12765_ _12629_/X _12765_/B VGND VGND VPWR VPWR _12766_/B sky130_fd_sc_hd__or2_4
XANTENNA__22885__B1 _21562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _21752_/A _14517_/B VGND VGND VPWR VPWR _14504_/Y sky130_fd_sc_hd__nand2_4
XPHY_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11716_/A VGND VGND VPWR VPWR _11717_/A sky130_fd_sc_hd__inv_2
X_18272_ _18205_/D _18272_/B VGND VGND VPWR VPWR _18273_/B sky130_fd_sc_hd__or2_4
XPHY_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ HWDATA[23] VGND VGND VPWR VPWR _15484_/X sky130_fd_sc_hd__buf_2
XPHY_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _13007_/B _12692_/Y _12695_/X VGND VGND VPWR VPWR _12696_/X sky130_fd_sc_hd__or3_4
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17223_ _17219_/Y _17222_/Y _16556_/X _17222_/Y VGND VGND VPWR VPWR _17223_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13378__B1 _11636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14435_ _15435_/A _14435_/B _14369_/B _14435_/D VGND VGND VPWR VPWR _14436_/B sky130_fd_sc_hd__and4_4
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ _11871_/A _11871_/B _25167_/Q VGND VGND VPWR VPWR _11647_/X sky130_fd_sc_hd__and3_4
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17154_ _17154_/A VGND VGND VPWR VPWR _17154_/Y sky130_fd_sc_hd__inv_2
X_14366_ _14366_/A VGND VGND VPWR VPWR _14366_/X sky130_fd_sc_hd__buf_2
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11578_ _11575_/Y _11569_/X _11576_/X _11577_/X VGND VGND VPWR VPWR _25206_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_92_0_HCLK clkbuf_8_93_0_HCLK/A VGND VGND VPWR VPWR _23668_/CLK sky130_fd_sc_hd__clkbuf_1
X_16105_ _16084_/A VGND VGND VPWR VPWR _16105_/X sky130_fd_sc_hd__buf_2
X_13317_ _13221_/A _13315_/X _13317_/C VGND VGND VPWR VPWR _13318_/C sky130_fd_sc_hd__and3_4
X_17085_ _17085_/A VGND VGND VPWR VPWR _24051_/D sky130_fd_sc_hd__inv_2
X_14297_ _14297_/A VGND VGND VPWR VPWR _14297_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23645__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16036_ _21257_/A _16035_/X _13480_/A VGND VGND VPWR VPWR _16036_/Y sky130_fd_sc_hd__a21oi_4
X_13248_ _13092_/A _19385_/A VGND VGND VPWR VPWR _13248_/X sky130_fd_sc_hd__or2_4
XFILLER_87_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16619__A1 _15657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13179_ _13278_/A _13177_/X _13178_/X VGND VGND VPWR VPWR _13179_/X sky130_fd_sc_hd__and3_4
XFILLER_69_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12092__A2_N _24545_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17987_ _17987_/A VGND VGND VPWR VPWR _17987_/X sky130_fd_sc_hd__buf_2
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19726_ _19726_/A VGND VGND VPWR VPWR _21325_/B sky130_fd_sc_hd__inv_2
XANTENNA__17562__A _17558_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16938_ _16936_/A _16938_/B _16937_/Y VGND VGND VPWR VPWR _24066_/D sky130_fd_sc_hd__and3_4
XFILLER_65_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19657_ _19656_/Y _19652_/X _19610_/X _19652_/X VGND VGND VPWR VPWR _23258_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11864__B1 _11708_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16869_ _16858_/A _16864_/Y _16868_/X VGND VGND VPWR VPWR _16869_/X sky130_fd_sc_hd__or3_4
XANTENNA__15055__B1 _15027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18608_ _23629_/Q _18608_/B VGND VGND VPWR VPWR _20279_/A sky130_fd_sc_hd__or2_4
X_19588_ _19575_/Y VGND VGND VPWR VPWR _19588_/X sky130_fd_sc_hd__buf_2
XFILLER_111_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24433__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21812__A _20966_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18539_ _18536_/A _18536_/B VGND VGND VPWR VPWR _18539_/Y sky130_fd_sc_hd__nand2_4
XFILLER_94_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19741__B1 _19714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21550_ _20235_/D _14016_/X _24812_/Q _21107_/X VGND VGND VPWR VPWR _21550_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13369__B1 _11616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20501_ _20484_/X _20500_/X _15357_/A _20488_/X VGND VGND VPWR VPWR _23713_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21481_ _21158_/A _19698_/Y VGND VGND VPWR VPWR _21481_/X sky130_fd_sc_hd__or2_4
XFILLER_119_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20432_ _20431_/X VGND VGND VPWR VPWR _23698_/D sky130_fd_sc_hd__inv_2
XANTENNA__13330__A _11643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23220_ _23292_/CLK _19766_/X VGND VGND VPWR VPWR _19764_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_119_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20363_ _23671_/Q _17174_/X VGND VGND VPWR VPWR _20363_/Y sky130_fd_sc_hd__nand2_4
XFILLER_31_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23151_ _25052_/CLK _23151_/D VGND VGND VPWR VPWR _23151_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_5_0_0_HCLK clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22102_ _20972_/A _19234_/Y VGND VGND VPWR VPWR _22102_/X sky130_fd_sc_hd__or2_4
XANTENNA__15530__A1 _15421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23082_ _23109_/CLK _23082_/D VGND VGND VPWR VPWR _23082_/Q sky130_fd_sc_hd__dfxtp_4
X_20294_ _14230_/Y _20273_/X _20287_/X _20293_/X VGND VGND VPWR VPWR _20295_/A sky130_fd_sc_hd__a211o_4
XANTENNA__25221__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22033_ _22032_/X VGND VGND VPWR VPWR _22033_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23628__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17283__B2 _17415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21706__B _21602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23984_ _23986_/CLK _23984_/D HRESETn VGND VGND VPWR VPWR _17239_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_25_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21906__A2 _21896_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22935_ _21864_/X _22933_/X _22530_/X _22934_/X VGND VGND VPWR VPWR _22935_/X sky130_fd_sc_hd__o22a_4
XANTENNA_clkbuf_3_7_0_HCLK_A clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19980__B1 _19455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16794__B1 _24416_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22866_ _16320_/A _16134_/X _21694_/X _22865_/X VGND VGND VPWR VPWR _22867_/C sky130_fd_sc_hd__a211o_4
XANTENNA__24174__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24605_ _24606_/CLK _24605_/D HRESETn VGND VGND VPWR VPWR _24605_/Q sky130_fd_sc_hd__dfrtp_4
X_21817_ _20962_/A _21815_/X _21816_/X VGND VGND VPWR VPWR _21817_/X sky130_fd_sc_hd__and3_4
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24103__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22797_ _15821_/X _22795_/X _22178_/A _22796_/X VGND VGND VPWR VPWR _22797_/X sky130_fd_sc_hd__o22a_4
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12550_ _12549_/Y VGND VGND VPWR VPWR _12550_/X sky130_fd_sc_hd__buf_2
XFILLER_24_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24536_ _25061_/CLK _15560_/X HRESETn VGND VGND VPWR VPWR _24536_/Q sky130_fd_sc_hd__dfrtp_4
X_21748_ _21747_/X VGND VGND VPWR VPWR _21748_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11501_ _11500_/X VGND VGND VPWR VPWR _11501_/X sky130_fd_sc_hd__buf_2
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12481_ _12478_/B VGND VGND VPWR VPWR _12481_/Y sky130_fd_sc_hd__inv_2
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24467_ _24042_/CLK _15711_/X HRESETn VGND VGND VPWR VPWR _20808_/A sky130_fd_sc_hd__dfrtp_4
X_21679_ _21675_/X _21678_/X _14486_/X VGND VGND VPWR VPWR _21688_/B sky130_fd_sc_hd__o21a_4
XFILLER_138_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ _20336_/A VGND VGND VPWR VPWR _20332_/A sky130_fd_sc_hd__inv_2
Xclkbuf_7_16_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_33_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12032__B1 _25144_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23418_ _23419_/CLK _23418_/D VGND VGND VPWR VPWR _17855_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24398_ _24399_/CLK _15903_/X HRESETn VGND VGND VPWR VPWR _24398_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_79_0_HCLK clkbuf_7_78_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_79_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14151_ _24838_/Q _14150_/X _14147_/A VGND VGND VPWR VPWR _14151_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_98_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17647__A _21153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23349_ _23350_/CLK _23349_/D VGND VGND VPWR VPWR _13106_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_137_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22272__B _21357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13102_ _13299_/A VGND VGND VPWR VPWR _13102_/X sky130_fd_sc_hd__buf_2
X_14082_ _14081_/Y _14079_/X _13665_/X _14079_/X VGND VGND VPWR VPWR _14082_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13033_ _13049_/A _23326_/Q VGND VGND VPWR VPWR _13033_/X sky130_fd_sc_hd__or2_4
X_17910_ _17878_/A _23440_/Q VGND VGND VPWR VPWR _17911_/C sky130_fd_sc_hd__or2_4
X_25019_ _25021_/CLK _25019_/D HRESETn VGND VGND VPWR VPWR _22419_/A sky130_fd_sc_hd__dfrtp_4
X_18890_ _23529_/Q VGND VGND VPWR VPWR _18890_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17841_ _17969_/A _17835_/X _17840_/X VGND VGND VPWR VPWR _17842_/C sky130_fd_sc_hd__or3_4
XFILLER_117_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20801__A _20800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24944__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14984_ _14984_/A VGND VGND VPWR VPWR _14984_/X sky130_fd_sc_hd__buf_2
X_17772_ _17878_/A _17772_/B VGND VGND VPWR VPWR _17772_/X sky130_fd_sc_hd__or2_4
XFILLER_66_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19511_ _19510_/Y VGND VGND VPWR VPWR _19511_/X sky130_fd_sc_hd__buf_2
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13935_ _13935_/A VGND VGND VPWR VPWR _13936_/A sky130_fd_sc_hd__buf_2
X_16723_ _21044_/A _17614_/A _24365_/Q _21839_/A VGND VGND VPWR VPWR _16726_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19971__B1 _19442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16654_ _16652_/X _16653_/X _11585_/A _24107_/Q _16647_/X VGND VGND VPWR VPWR _16654_/X
+ sky130_fd_sc_hd__a32o_4
X_19442_ _19442_/A VGND VGND VPWR VPWR _19442_/X sky130_fd_sc_hd__buf_2
X_13866_ _13866_/A _13866_/B VGND VGND VPWR VPWR _13866_/Y sky130_fd_sc_hd__nand2_4
XFILLER_62_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15605_ _12559_/Y _15604_/X _15350_/X _15604_/X VGND VGND VPWR VPWR _24523_/D sky130_fd_sc_hd__a2bb2o_4
X_12817_ _22203_/A _22187_/A _12815_/Y _12816_/Y VGND VGND VPWR VPWR _12821_/C sky130_fd_sc_hd__o22a_4
X_16585_ _16583_/Y _16584_/X _16254_/X _16584_/X VGND VGND VPWR VPWR _16585_/X sky130_fd_sc_hd__a2bb2o_4
X_19373_ _19372_/Y VGND VGND VPWR VPWR _19373_/X sky130_fd_sc_hd__buf_2
X_13797_ _13797_/A _14073_/B _13797_/C _13789_/Y VGND VGND VPWR VPWR _13798_/A sky130_fd_sc_hd__or4_4
XFILLER_50_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21125__A3 _21432_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15536_ _15535_/X VGND VGND VPWR VPWR _15558_/A sky130_fd_sc_hd__buf_2
X_18324_ _18214_/Y _18301_/B _18322_/B _18237_/X VGND VGND VPWR VPWR _18325_/A sky130_fd_sc_hd__a211o_4
X_12748_ _12581_/Y _12742_/B VGND VGND VPWR VPWR _12749_/C sky130_fd_sc_hd__nand2_4
XFILLER_37_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21530__B1 _21529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18255_ _18240_/X VGND VGND VPWR VPWR _18260_/B sky130_fd_sc_hd__inv_2
XANTENNA__23897__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15467_ _15368_/X _15461_/X _15320_/X _24576_/Q _15466_/X VGND VGND VPWR VPWR _24576_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_8_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12679_ _12550_/X _12571_/Y _12679_/C _12694_/B VGND VGND VPWR VPWR _12679_/X sky130_fd_sc_hd__or4_4
XFILLER_30_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17206_ _17213_/A VGND VGND VPWR VPWR _17206_/X sky130_fd_sc_hd__buf_2
X_14418_ _14378_/Y _14417_/X _14412_/X _14415_/X _14377_/A VGND VGND VPWR VPWR _14418_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23826__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18186_ _16119_/Y _18211_/A _16123_/A _18167_/Y VGND VGND VPWR VPWR _18190_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12023__B1 _12001_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15398_ _24587_/Q VGND VGND VPWR VPWR _15398_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22463__A _22463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17137_ _24038_/Q _17137_/B VGND VGND VPWR VPWR _17139_/B sky130_fd_sc_hd__or2_4
X_14349_ _20271_/A VGND VGND VPWR VPWR _14349_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17068_ _17070_/B VGND VGND VPWR VPWR _17074_/B sky130_fd_sc_hd__inv_2
XANTENNA__21079__A _20852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16019_ _14434_/A _16014_/C VGND VGND VPWR VPWR _16019_/X sky130_fd_sc_hd__and2_4
XANTENNA__17265__A1 _25192_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21807__A _20833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24685__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15805__A _15439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24614__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19709_ _19709_/A VGND VGND VPWR VPWR _19709_/Y sky130_fd_sc_hd__inv_2
X_20981_ _20975_/X _20980_/X _20968_/X VGND VGND VPWR VPWR _20981_/X sky130_fd_sc_hd__o21a_4
XFILLER_66_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15028__B1 _15027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0_0_HCLK_A clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17014__A2_N _17021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13325__A _13324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22720_ _12619_/Y _20910_/X _12853_/Y _22029_/X VGND VGND VPWR VPWR _22720_/X sky130_fd_sc_hd__o22a_4
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21542__A _21848_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22849__B1 _24571_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22651_ _22651_/A _22651_/B VGND VGND VPWR VPWR _22651_/X sky130_fd_sc_hd__and2_4
XFILLER_34_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21602_ _21602_/A _21569_/X _21602_/C _21601_/Y VGND VGND VPWR VPWR _21602_/X sky130_fd_sc_hd__or4_4
XANTENNA__15540__A _19445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19012__A _19012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16528__B1 _16100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22582_ _16078_/A _22350_/X _22581_/X VGND VGND VPWR VPWR _22582_/X sky130_fd_sc_hd__o21a_4
XFILLER_90_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24321_ _24071_/CLK _24321_/D HRESETn VGND VGND VPWR VPWR _24321_/Q sky130_fd_sc_hd__dfrtp_4
X_21533_ _21400_/X _21532_/X _13419_/Y _21400_/X VGND VGND VPWR VPWR _21533_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18851__A _13039_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24252_ _24225_/CLK _24252_/D HRESETn VGND VGND VPWR VPWR _16310_/A sky130_fd_sc_hd__dfrtp_4
X_21464_ _21350_/A _21464_/B _21463_/X VGND VGND VPWR VPWR _21464_/X sky130_fd_sc_hd__and3_4
XANTENNA__22373__A _22373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23203_ _24008_/CLK _23203_/D VGND VGND VPWR VPWR _13170_/B sky130_fd_sc_hd__dfxtp_4
X_20415_ _20414_/X VGND VGND VPWR VPWR _20416_/A sky130_fd_sc_hd__buf_2
X_21395_ _21391_/X _21394_/X _21242_/X VGND VGND VPWR VPWR _21396_/C sky130_fd_sc_hd__o21a_4
X_24183_ _24113_/CLK _16494_/X HRESETn VGND VGND VPWR VPWR _16492_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_135_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23134_ _23992_/CLK _19992_/X VGND VGND VPWR VPWR _23134_/Q sky130_fd_sc_hd__dfxtp_4
X_20346_ _14059_/Y _20344_/X _20401_/A _20345_/X VGND VGND VPWR VPWR _20347_/A sky130_fd_sc_hd__a211o_4
X_20277_ _23629_/Q _18608_/B VGND VGND VPWR VPWR _20279_/B sky130_fd_sc_hd__nand2_4
XFILLER_122_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23065_ _23664_/CLK scl_oen_o_S5 VGND VGND VPWR VPWR _20720_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__11915__A1_N _11913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12404__A _21104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17256__A1 _25214_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22016_ _21719_/A _22014_/X _16368_/Y _22015_/X VGND VGND VPWR VPWR _22016_/X sky130_fd_sc_hd__o22a_4
XFILLER_7_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20621__A _20647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24355__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22001__B2 _21051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11981_ _13398_/A VGND VGND VPWR VPWR _11981_/X sky130_fd_sc_hd__buf_2
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23967_ _24378_/CLK _23967_/D HRESETn VGND VGND VPWR VPWR _17482_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19150__A2_N _19146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13720_ _13754_/A _13742_/C _13770_/A _13780_/B VGND VGND VPWR VPWR _13720_/X sky130_fd_sc_hd__or4_4
XFILLER_95_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22552__A2 _21896_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22918_ _21546_/X _22915_/Y _22423_/X _22917_/X VGND VGND VPWR VPWR _22918_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21416__A1_N _21040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23898_ _23898_/CLK _18062_/Y HRESETn VGND VGND VPWR VPWR _21491_/A sky130_fd_sc_hd__dfstp_4
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22548__A _22548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13651_ _22449_/A _13649_/X _11585_/X _13649_/X VGND VGND VPWR VPWR _24939_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22849_ _23020_/B _22848_/X _22839_/X _24571_/Q _20833_/X VGND VGND VPWR VPWR _22849_/X
+ sky130_fd_sc_hd__a32o_4
X_12602_ _12594_/X _12597_/X _12599_/X _12601_/X VGND VGND VPWR VPWR _12632_/A sky130_fd_sc_hd__or4_4
XANTENNA__22267__B _22314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16370_ _16368_/Y _16364_/X _16369_/X _16364_/X VGND VGND VPWR VPWR _24229_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13582_ _13564_/X _13580_/X _13581_/Y _13576_/X _24958_/Q VGND VGND VPWR VPWR _24958_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16519__B1 _16087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15321_ _13358_/X VGND VGND VPWR VPWR _15322_/A sky130_fd_sc_hd__buf_2
XFILLER_12_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23990__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12533_ _12389_/X _12535_/B _12532_/Y VGND VGND VPWR VPWR _25073_/D sky130_fd_sc_hd__o21a_4
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24519_ _24523_/CLK _24519_/D HRESETn VGND VGND VPWR VPWR _24519_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18040_ _18020_/X _18039_/X _18020_/X _18039_/X VGND VGND VPWR VPWR _18040_/X sky130_fd_sc_hd__a2bb2o_4
X_15252_ _15250_/X _23765_/Q _15251_/Y _13761_/A _15245_/X VGND VGND VPWR VPWR _15252_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12005__B1 _11631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12464_ _12498_/A _12495_/A _12502_/A _12409_/X VGND VGND VPWR VPWR _12464_/X sky130_fd_sc_hd__or4_4
XANTENNA__15742__A1 _15421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25143__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14203_ _20193_/A _14200_/X _13663_/X _14202_/X VGND VGND VPWR VPWR _14203_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15183_ _15165_/A _15183_/B _15183_/C VGND VGND VPWR VPWR _15183_/X sky130_fd_sc_hd__and3_4
X_12395_ _12408_/C _24473_/Q _12389_/X _24470_/Q VGND VGND VPWR VPWR _12395_/X sky130_fd_sc_hd__a2bb2o_4
X_14134_ _14126_/X _14133_/X _24992_/Q _14131_/X VGND VGND VPWR VPWR _24846_/D sky130_fd_sc_hd__o22a_4
X_19991_ _19990_/Y VGND VGND VPWR VPWR _19991_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_103_0_HCLK clkbuf_7_51_0_HCLK/X VGND VGND VPWR VPWR _24017_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_4_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14065_ _14064_/Y _14060_/X _13645_/X _14048_/A VGND VGND VPWR VPWR _14065_/X sky130_fd_sc_hd__a2bb2o_4
X_18942_ _17685_/B VGND VGND VPWR VPWR _18942_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_166_0_HCLK clkbuf_7_83_0_HCLK/X VGND VGND VPWR VPWR _24740_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_9_0_HCLK clkbuf_6_4_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13016_ _13016_/A VGND VGND VPWR VPWR _13042_/A sky130_fd_sc_hd__buf_2
X_18873_ _24732_/Q _18873_/B _13461_/X VGND VGND VPWR VPWR _18873_/X sky130_fd_sc_hd__or3_4
X_17824_ _17955_/A _17815_/X _17824_/C VGND VGND VPWR VPWR _17824_/X sky130_fd_sc_hd__and3_4
XANTENNA__24096__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14967_ _14966_/Y _24285_/Q _14966_/Y _24285_/Q VGND VGND VPWR VPWR _14972_/B sky130_fd_sc_hd__a2bb2o_4
X_17755_ _17927_/A _23533_/Q VGND VGND VPWR VPWR _17755_/X sky130_fd_sc_hd__or2_4
XFILLER_130_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13145__A _13169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16706_ _24367_/Q _16704_/A _15984_/Y _17595_/C VGND VGND VPWR VPWR _16707_/D sky130_fd_sc_hd__o22a_4
X_13918_ _13891_/A VGND VGND VPWR VPWR _20179_/C sky130_fd_sc_hd__buf_2
XANTENNA__19748__A2_N _19743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14898_ _24676_/Q VGND VGND VPWR VPWR _14898_/Y sky130_fd_sc_hd__inv_2
X_17686_ _17702_/A _17684_/X _17685_/X VGND VGND VPWR VPWR _17686_/X sky130_fd_sc_hd__and3_4
XANTENNA__16993__A1_N _24306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19425_ _19417_/Y VGND VGND VPWR VPWR _19425_/X sky130_fd_sc_hd__buf_2
X_13849_ _13830_/C VGND VGND VPWR VPWR _13849_/Y sky130_fd_sc_hd__inv_2
X_16637_ _16624_/X _16625_/X HWDATA[23] _24116_/Q _16622_/X VGND VGND VPWR VPWR _16637_/X
+ sky130_fd_sc_hd__a32o_4
X_19356_ _19354_/Y _19350_/X _19311_/X _19355_/X VGND VGND VPWR VPWR _19356_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21892__A2_N _20818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16568_ _16566_/A VGND VGND VPWR VPWR _16575_/A sky130_fd_sc_hd__inv_2
XFILLER_128_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18307_ _18213_/D _18307_/B VGND VGND VPWR VPWR _18311_/B sky130_fd_sc_hd__or2_4
X_15519_ _12125_/Y _15518_/X _15393_/X _15518_/X VGND VGND VPWR VPWR _24550_/D sky130_fd_sc_hd__a2bb2o_4
X_16499_ _16499_/A VGND VGND VPWR VPWR _16499_/X sky130_fd_sc_hd__buf_2
X_19287_ _21928_/B _19284_/X _11839_/X _19284_/X VGND VGND VPWR VPWR _23389_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23660__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18238_ _18179_/Y _18231_/X _18237_/X _18234_/B VGND VGND VPWR VPWR _18239_/A sky130_fd_sc_hd__a211o_4
XANTENNA__12000__A1_N _11999_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18169_ _16123_/A _18167_/Y _24329_/Q _18216_/A VGND VGND VPWR VPWR _18172_/B sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_62_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_62_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20200_ _20200_/A VGND VGND VPWR VPWR _20200_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16289__A2 _16276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21180_ _21400_/A VGND VGND VPWR VPWR _21180_/X sky130_fd_sc_hd__buf_2
XANTENNA__18683__B1 _16671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20131_ _20131_/A VGND VGND VPWR VPWR _20131_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20062_ _20062_/A VGND VGND VPWR VPWR _20062_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17238__B2 _25221_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13039__B _13039_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15535__A _14369_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24870_ _24870_/CLK _14051_/X HRESETn VGND VGND VPWR VPWR _14050_/A sky130_fd_sc_hd__dfstp_4
XFILLER_100_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23821_ _23826_/CLK _23821_/D HRESETn VGND VGND VPWR VPWR _23821_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19935__B1 _19452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13055__A _13054_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23752_ _24180_/CLK _23752_/D HRESETn VGND VGND VPWR VPWR _23752_/Q sky130_fd_sc_hd__dfrtp_4
X_20964_ _20964_/A _20964_/B VGND VGND VPWR VPWR _20967_/B sky130_fd_sc_hd__or2_4
XFILLER_54_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22703_ _22703_/A _22703_/B VGND VGND VPWR VPWR _22703_/X sky130_fd_sc_hd__or2_4
XFILLER_14_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23683_ _24769_/CLK sda_i_S5 HRESETn VGND VGND VPWR VPWR _23684_/D sky130_fd_sc_hd__dfrtp_4
X_20895_ _20894_/X VGND VGND VPWR VPWR _20896_/D sky130_fd_sc_hd__inv_2
XFILLER_110_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23748__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22634_ _22629_/A VGND VGND VPWR VPWR _22634_/X sky130_fd_sc_hd__buf_2
XFILLER_10_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22565_ _22565_/A _15655_/A VGND VGND VPWR VPWR _22565_/X sky130_fd_sc_hd__and2_4
XFILLER_10_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24304_ _24037_/CLK _24304_/D HRESETn VGND VGND VPWR VPWR _16181_/A sky130_fd_sc_hd__dfrtp_4
X_21516_ _14529_/X VGND VGND VPWR VPWR _21519_/A sky130_fd_sc_hd__buf_2
X_22496_ _22472_/X _22476_/X _22482_/Y _22495_/X VGND VGND VPWR VPWR HRDATA[15] sky130_fd_sc_hd__a211o_4
XFILLER_108_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17197__A _13619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24235_ _23840_/CLK _16355_/X HRESETn VGND VGND VPWR VPWR _16354_/A sky130_fd_sc_hd__dfrtp_4
X_21447_ _21447_/A _21446_/X VGND VGND VPWR VPWR _21457_/C sky130_fd_sc_hd__and2_4
X_12180_ _12180_/A _12180_/B _12265_/C _12091_/Y VGND VGND VPWR VPWR _12180_/X sky130_fd_sc_hd__or4_4
XANTENNA__11957__B _11956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18674__B1 _17205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24166_ _24167_/CLK _16536_/X HRESETn VGND VGND VPWR VPWR _16534_/A sky130_fd_sc_hd__dfrtp_4
X_21378_ _21378_/A _19853_/Y VGND VGND VPWR VPWR _21379_/C sky130_fd_sc_hd__or2_4
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15488__B1 _15350_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23117_ _23388_/CLK _20037_/X VGND VGND VPWR VPWR _20033_/A sky130_fd_sc_hd__dfxtp_4
X_20329_ _14247_/Y _18624_/A _18607_/A _18620_/Y VGND VGND VPWR VPWR _20330_/B sky130_fd_sc_hd__o22a_4
XFILLER_134_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24097_ _24094_/CLK _24097_/D HRESETn VGND VGND VPWR VPWR _24097_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24536__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_239_0_HCLK clkbuf_8_239_0_HCLK/A VGND VGND VPWR VPWR _24180_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21025__A2 _20988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23048_ VGND VGND VPWR VPWR _23048_/HI scl_o_S4 sky130_fd_sc_hd__conb_1
XFILLER_89_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15870_ _24410_/Q VGND VGND VPWR VPWR _15870_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14821_ _14821_/A VGND VGND VPWR VPWR _14821_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24999_ _24998_/CLK _24999_/D HRESETn VGND VGND VPWR VPWR _24999_/Q sky130_fd_sc_hd__dfrtp_4
X_14752_ _24687_/Q VGND VGND VPWR VPWR _14869_/B sky130_fd_sc_hd__inv_2
X_17540_ _17539_/X VGND VGND VPWR VPWR _23966_/D sky130_fd_sc_hd__inv_2
X_11964_ _11964_/A VGND VGND VPWR VPWR _22982_/A sky130_fd_sc_hd__buf_2
XFILLER_44_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13703_ _13697_/X _13702_/X _24858_/Q _13693_/X VGND VGND VPWR VPWR _13703_/X sky130_fd_sc_hd__o22a_4
X_17471_ _17463_/X _17470_/Y _23976_/Q _17462_/Y VGND VGND VPWR VPWR _17471_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14683_ _14683_/A _14682_/X VGND VGND VPWR VPWR _14683_/Y sky130_fd_sc_hd__nor2_4
X_11895_ _23785_/Q _11882_/B _11894_/Y VGND VGND VPWR VPWR _20688_/A sky130_fd_sc_hd__o21a_4
X_19210_ _19209_/Y _19204_/X _19120_/X _19196_/A VGND VGND VPWR VPWR _23415_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13634_ _24944_/Q VGND VGND VPWR VPWR _13634_/Y sky130_fd_sc_hd__inv_2
X_16422_ _16420_/Y _16421_/X _16334_/X _16421_/X VGND VGND VPWR VPWR _24211_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16353_ _16351_/Y _16347_/X _15369_/X _16352_/X VGND VGND VPWR VPWR _24236_/D sky130_fd_sc_hd__a2bb2o_4
X_19141_ _23439_/Q VGND VGND VPWR VPWR _19141_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12777__B2 _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13565_ _13564_/X VGND VGND VPWR VPWR _13566_/B sky130_fd_sc_hd__inv_2
XANTENNA__16730__A2_N _22473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15304_ _15300_/Y VGND VGND VPWR VPWR _15304_/X sky130_fd_sc_hd__buf_2
X_12516_ _12345_/X _12515_/X _12427_/X VGND VGND VPWR VPWR _12516_/Y sky130_fd_sc_hd__a21oi_4
X_19072_ _19070_/Y _19071_/X _18959_/X _19071_/X VGND VGND VPWR VPWR _23465_/D sky130_fd_sc_hd__a2bb2o_4
X_16284_ _14916_/Y _16282_/X _15890_/X _16282_/X VGND VGND VPWR VPWR _16284_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13496_ _20499_/A _20499_/B _20499_/C _22656_/A VGND VGND VPWR VPWR _13497_/D sky130_fd_sc_hd__or4_4
XFILLER_12_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15235_ _15234_/X VGND VGND VPWR VPWR _15235_/Y sky130_fd_sc_hd__inv_2
X_18023_ _18023_/A VGND VGND VPWR VPWR _18023_/X sky130_fd_sc_hd__buf_2
X_12447_ _12415_/A _12458_/A VGND VGND VPWR VPWR _12448_/B sky130_fd_sc_hd__or2_4
Xclkbuf_6_49_0_HCLK clkbuf_6_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_99_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15166_ _15161_/A _15161_/B _15126_/X _15163_/B VGND VGND VPWR VPWR _15166_/X sky130_fd_sc_hd__a211o_4
X_12378_ _12415_/B _22736_/A _25080_/Q _12316_/Y VGND VGND VPWR VPWR _12387_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22461__B2 _22460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14117_ _14107_/Y _14116_/X _13488_/X VGND VGND VPWR VPWR _14117_/Y sky130_fd_sc_hd__a21oi_4
X_15097_ _14867_/A _15085_/X _15097_/C VGND VGND VPWR VPWR _15097_/X sky130_fd_sc_hd__and3_4
X_19974_ _23140_/Q VGND VGND VPWR VPWR _21777_/B sky130_fd_sc_hd__inv_2
XFILLER_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24277__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14048_ _14048_/A VGND VGND VPWR VPWR _14048_/X sky130_fd_sc_hd__buf_2
X_18925_ _18924_/Y _18922_/X _18880_/X _18922_/X VGND VGND VPWR VPWR _23517_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22213__A1 _21870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21357__A _21357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24206__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18856_ _13063_/B VGND VGND VPWR VPWR _18856_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19090__B1 _19089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17807_ _17916_/A _17807_/B VGND VGND VPWR VPWR _17809_/B sky130_fd_sc_hd__or2_4
XFILLER_55_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17640__A1 _17639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_4_0_HCLK clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_4_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18787_ _17745_/B VGND VGND VPWR VPWR _18787_/Y sky130_fd_sc_hd__inv_2
X_15999_ _21044_/A VGND VGND VPWR VPWR _15999_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17738_ _17738_/A _17738_/B _17737_/X VGND VGND VPWR VPWR _17739_/C sky130_fd_sc_hd__or3_4
XFILLER_63_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22188__A _20866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21092__A _20861_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19393__B2 _19372_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17669_ _13406_/B _17656_/Y _17665_/X VGND VGND VPWR VPWR _17669_/X sky130_fd_sc_hd__o21a_4
XFILLER_90_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15090__A _15087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19408_ _13249_/B VGND VGND VPWR VPWR _19408_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23841__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12217__B1 _12195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20680_ _20676_/X VGND VGND VPWR VPWR _20680_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25065__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22916__A _24495_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19339_ _19338_/Y _19334_/X _19201_/X _19334_/X VGND VGND VPWR VPWR _19339_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22350_ _22616_/A VGND VGND VPWR VPWR _22350_/X sky130_fd_sc_hd__buf_2
XANTENNA__14509__A2 _14484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21301_ _14818_/A _20931_/X _21299_/X _21300_/Y VGND VGND VPWR VPWR _21302_/C sky130_fd_sc_hd__a211o_4
X_22281_ _20900_/A VGND VGND VPWR VPWR _22281_/X sky130_fd_sc_hd__buf_2
XANTENNA__17448__C _21363_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24020_ _24643_/CLK _17195_/X HRESETn VGND VGND VPWR VPWR _20733_/A sky130_fd_sc_hd__dfrtp_4
X_21232_ _21224_/X _21230_/X _21231_/X VGND VGND VPWR VPWR _21244_/B sky130_fd_sc_hd__o21a_4
XFILLER_116_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16255__A1_N _14960_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21163_ _17644_/A VGND VGND VPWR VPWR _21350_/A sky130_fd_sc_hd__buf_2
XANTENNA__11668__A2_N _22450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22528__A2_N _22259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20114_ _20114_/A VGND VGND VPWR VPWR _20982_/B sky130_fd_sc_hd__inv_2
XFILLER_28_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15485__A3 _15484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21094_ _21275_/A _21093_/X _16616_/Y _20863_/A VGND VGND VPWR VPWR _21094_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22204__B2 _22167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20045_ _23113_/Q VGND VGND VPWR VPWR _21475_/B sky130_fd_sc_hd__inv_2
X_24922_ _24879_/CLK _13691_/X HRESETn VGND VGND VPWR VPWR _20201_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_63_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_69_0_HCLK clkbuf_8_69_0_HCLK/A VGND VGND VPWR VPWR _23641_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24853_ _24980_/CLK _14106_/X HRESETn VGND VGND VPWR VPWR _24853_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12401__B _12401_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17480__A _22853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23929__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23804_ _24017_/CLK _18634_/X HRESETn VGND VGND VPWR VPWR _20717_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_38_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24784_ _24788_/CLK _24784_/D HRESETn VGND VGND VPWR VPWR _14306_/A sky130_fd_sc_hd__dfrtp_4
X_21996_ _15322_/A _21993_/X _21994_/X _11614_/A _21995_/X VGND VGND VPWR VPWR _21996_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_73_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23735_ _24167_/CLK _23735_/D HRESETn VGND VGND VPWR VPWR _20590_/A sky130_fd_sc_hd__dfrtp_4
X_20947_ _20946_/X _20947_/B VGND VGND VPWR VPWR _20947_/X sky130_fd_sc_hd__or2_4
XPHY_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16096__A _16096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _23918_/Q VGND VGND VPWR VPWR _11680_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14748__A2 _14747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23666_ _23661_/CLK _23666_/D HRESETn VGND VGND VPWR VPWR _23666_/Q sky130_fd_sc_hd__dfstp_4
X_20878_ _21072_/A _20878_/B VGND VGND VPWR VPWR _20878_/Y sky130_fd_sc_hd__nor2_4
XPHY_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22617_ _24274_/Q _22616_/X _22338_/X VGND VGND VPWR VPWR _22617_/X sky130_fd_sc_hd__o21a_4
XFILLER_35_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22140__B1 _21581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23597_ _25009_/CLK _18695_/X VGND VGND VPWR VPWR _23597_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13350_ _13350_/A VGND VGND VPWR VPWR _13350_/Y sky130_fd_sc_hd__inv_2
X_22548_ _22548_/A VGND VGND VPWR VPWR _22549_/A sky130_fd_sc_hd__buf_2
X_12301_ _12091_/Y _12192_/B _12203_/X _12299_/B VGND VGND VPWR VPWR _12302_/A sky130_fd_sc_hd__a211o_4
XANTENNA__13708__B1 _23126_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24788__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13281_ _13146_/A _19411_/A VGND VGND VPWR VPWR _13281_/X sky130_fd_sc_hd__or2_4
X_22479_ _22479_/A _22265_/B VGND VGND VPWR VPWR _22479_/X sky130_fd_sc_hd__and2_4
XFILLER_5_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15020_ _15045_/A _15042_/A _15019_/X VGND VGND VPWR VPWR _15020_/X sky130_fd_sc_hd__or3_4
XANTENNA__24717__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12232_ _12172_/A _12232_/B VGND VGND VPWR VPWR _12234_/B sky130_fd_sc_hd__or2_4
X_24218_ _24192_/CLK _24218_/D HRESETn VGND VGND VPWR VPWR _24218_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22653__A1_N _12412_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25198_ _23957_/CLK _25198_/D HRESETn VGND VGND VPWR VPWR _25198_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_5_3_0_HCLK_A clkbuf_5_2_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12163_ _12502_/A VGND VGND VPWR VPWR _12423_/A sky130_fd_sc_hd__buf_2
XFILLER_68_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24149_ _24098_/CLK _24149_/D HRESETn VGND VGND VPWR VPWR _24149_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24370__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21177__A _20753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12094_ _25121_/Q VGND VGND VPWR VPWR _12094_/Y sky130_fd_sc_hd__inv_2
X_16971_ _16218_/Y _17031_/A _16218_/Y _17031_/A VGND VGND VPWR VPWR _16972_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18710_ _23591_/Q VGND VGND VPWR VPWR _18710_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15881__B1 _11598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15922_ _15921_/X VGND VGND VPWR VPWR _15922_/X sky130_fd_sc_hd__buf_2
XANTENNA__19072__B1 _18959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19690_ _19686_/Y _19689_/X _19597_/X _19689_/X VGND VGND VPWR VPWR _23246_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18641_ _19779_/B VGND VGND VPWR VPWR _19862_/B sky130_fd_sc_hd__buf_2
X_15853_ _24416_/Q VGND VGND VPWR VPWR _15853_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15633__B1 _15286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14804_ _14882_/A _24153_/Q _14882_/A _24153_/Q VGND VGND VPWR VPWR _14804_/X sky130_fd_sc_hd__a2bb2o_4
X_18572_ _16345_/A _23829_/Q _16345_/Y _18434_/D VGND VGND VPWR VPWR _18576_/A sky130_fd_sc_hd__o22a_4
X_12996_ _12972_/A _12972_/B _12922_/A _12993_/Y VGND VGND VPWR VPWR _12996_/X sky130_fd_sc_hd__a211o_4
X_15784_ _15781_/X _15763_/X _16093_/A _22385_/A _15779_/X VGND VGND VPWR VPWR _24442_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_45_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17523_ _17505_/C _17515_/B VGND VGND VPWR VPWR _17524_/A sky130_fd_sc_hd__or2_4
X_11947_ _15414_/A VGND VGND VPWR VPWR _16301_/A sky130_fd_sc_hd__buf_2
X_14735_ _24701_/Q VGND VGND VPWR VPWR _14876_/C sky130_fd_sc_hd__inv_2
XFILLER_75_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14666_ _14657_/X _14665_/Y _14045_/A _14657_/X VGND VGND VPWR VPWR _14666_/X sky130_fd_sc_hd__a2bb2o_4
X_17454_ _17451_/Y _17453_/X _23976_/Q _17452_/A VGND VGND VPWR VPWR _17454_/X sky130_fd_sc_hd__o22a_4
X_11878_ _11871_/B _11867_/X _11877_/Y VGND VGND VPWR VPWR _25165_/D sky130_fd_sc_hd__o21a_4
X_13617_ _22439_/B VGND VGND VPWR VPWR _13618_/A sky130_fd_sc_hd__buf_2
X_16405_ _16404_/Y _16402_/X _11536_/X _16402_/X VGND VGND VPWR VPWR _24218_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_12_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_12_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_14597_ _19189_/B _14587_/X _14592_/B VGND VGND VPWR VPWR _14597_/X sky130_fd_sc_hd__a21o_4
X_17385_ _17382_/C _17382_/D VGND VGND VPWR VPWR _17386_/B sky130_fd_sc_hd__or2_4
XANTENNA__22131__B1 _24552_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19124_ _19123_/X VGND VGND VPWR VPWR _19137_/A sky130_fd_sc_hd__inv_2
X_13548_ _20883_/A _20881_/A _24965_/Q VGND VGND VPWR VPWR _24963_/D sky130_fd_sc_hd__a21o_4
X_16336_ _24242_/Q VGND VGND VPWR VPWR _16336_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22682__B2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12383__A2_N _24493_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16267_ _14933_/Y _16262_/X _16266_/X _16262_/X VGND VGND VPWR VPWR _16267_/X sky130_fd_sc_hd__a2bb2o_4
X_19055_ _23470_/Q VGND VGND VPWR VPWR _19055_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13479_ _21700_/A _13478_/Y _13402_/A _13478_/A VGND VGND VPWR VPWR _13479_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16684__A2_N _23012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24458__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15218_ _15218_/A _15218_/B VGND VGND VPWR VPWR _15219_/B sky130_fd_sc_hd__or2_4
X_18006_ _17979_/X _11944_/X VGND VGND VPWR VPWR _18007_/A sky130_fd_sc_hd__or2_4
X_16198_ _16198_/A VGND VGND VPWR VPWR _16198_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24025__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15149_ _15138_/A _15146_/X _15148_/Y VGND VGND VPWR VPWR _24675_/D sky130_fd_sc_hd__o21a_4
XFILLER_99_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22985__A2 _22505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15467__A3 _15320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19957_ _23146_/Q VGND VGND VPWR VPWR _19957_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24040__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_222_0_HCLK clkbuf_8_223_0_HCLK/A VGND VGND VPWR VPWR _24262_/CLK sky130_fd_sc_hd__clkbuf_1
X_18908_ _17834_/B VGND VGND VPWR VPWR _18908_/Y sky130_fd_sc_hd__inv_2
X_19888_ _21960_/B _19885_/X _19818_/X _19885_/X VGND VGND VPWR VPWR _19888_/X sky130_fd_sc_hd__a2bb2o_4
X_18839_ _18837_/Y _18833_/X _15550_/X _18838_/X VGND VGND VPWR VPWR _23548_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18810__B1 _18764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21850_ _21850_/A _21849_/X VGND VGND VPWR VPWR _21855_/C sky130_fd_sc_hd__and2_4
XFILLER_83_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20801_ _20800_/X VGND VGND VPWR VPWR _20801_/X sky130_fd_sc_hd__buf_2
XFILLER_93_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21781_ _21383_/A _21781_/B VGND VGND VPWR VPWR _21781_/X sky130_fd_sc_hd__or2_4
XANTENNA__13333__A _13333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23520_ _23560_/CLK _23520_/D VGND VGND VPWR VPWR _18915_/A sky130_fd_sc_hd__dfxtp_4
X_20732_ _23660_/Q _23661_/Q _20733_/B VGND VGND VPWR VPWR _23660_/D sky130_fd_sc_hd__o21a_4
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20920__A1 _20910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23451_ _23440_/CLK _23451_/D VGND VGND VPWR VPWR _17807_/B sky130_fd_sc_hd__dfxtp_4
X_20663_ _23752_/Q VGND VGND VPWR VPWR _20663_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22365__B _21979_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22402_ _22264_/X _22401_/X _16354_/Y _16305_/X VGND VGND VPWR VPWR _22402_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23382_ _23374_/CLK _23382_/D VGND VGND VPWR VPWR _13023_/B sky130_fd_sc_hd__dfxtp_4
X_20594_ _23736_/Q VGND VGND VPWR VPWR _20594_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24881__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20684__B1 _11708_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25121_ _25123_/CLK _12241_/X HRESETn VGND VGND VPWR VPWR _25121_/Q sky130_fd_sc_hd__dfrtp_4
X_22333_ _21570_/X VGND VGND VPWR VPWR _22334_/A sky130_fd_sc_hd__buf_2
XFILLER_109_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15155__A2 _15123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24199__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14363__B1 sda_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25052_ _25052_/CLK _25052_/D HRESETn VGND VGND VPWR VPWR _12609_/A sky130_fd_sc_hd__dfrtp_4
X_22264_ _22226_/A VGND VGND VPWR VPWR _22264_/X sky130_fd_sc_hd__buf_2
XFILLER_121_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24128__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24003_ _25217_/CLK _17360_/X HRESETn VGND VGND VPWR VPWR _17306_/A sky130_fd_sc_hd__dfrtp_4
X_21215_ _21378_/A _21215_/B VGND VGND VPWR VPWR _21215_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_32_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_32_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22195_ _20753_/A VGND VGND VPWR VPWR _22195_/X sky130_fd_sc_hd__buf_2
X_21146_ _21336_/A _21146_/B VGND VGND VPWR VPWR _21146_/X sky130_fd_sc_hd__or2_4
XANTENNA__13469__A2 _13480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22189__B1 _12582_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15863__B1 _15775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22728__A2 _21896_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19054__B1 _18964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21077_ _21073_/X _21074_/X _21075_/X _21076_/X VGND VGND VPWR VPWR _21077_/X sky130_fd_sc_hd__or4_4
XANTENNA__12412__A _12412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20028_ _21326_/B _20027_/X _19728_/X _20027_/X VGND VGND VPWR VPWR _20028_/X sky130_fd_sc_hd__a2bb2o_4
X_24905_ _24902_/CLK _13907_/X HRESETn VGND VGND VPWR VPWR _24905_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15615__B1 _24516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23763__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12850_ _12972_/A _15797_/A _22921_/A _12849_/Y VGND VGND VPWR VPWR _12856_/B sky130_fd_sc_hd__a2bb2o_4
X_24836_ _24851_/CLK _14156_/X HRESETn VGND VGND VPWR VPWR _12049_/A sky130_fd_sc_hd__dfrtp_4
X_11801_ _17448_/B RsRx_S1 VGND VGND VPWR VPWR _11801_/X sky130_fd_sc_hd__or2_4
XFILLER_132_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16762__A1_N _24416_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12781_ _22826_/A VGND VGND VPWR VPWR _12781_/Y sky130_fd_sc_hd__inv_2
X_24767_ _24968_/CLK _14391_/X HRESETn VGND VGND VPWR VPWR _24767_/Q sky130_fd_sc_hd__dfrtp_4
X_21979_ _21848_/B VGND VGND VPWR VPWR _21979_/X sky130_fd_sc_hd__buf_2
XFILLER_92_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14519_/Y _14507_/Y _21752_/A _14506_/X VGND VGND VPWR VPWR _14520_/X sky130_fd_sc_hd__o22a_4
XPHY_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11732_ _11732_/A _11732_/B VGND VGND VPWR VPWR _11733_/B sky130_fd_sc_hd__and2_4
XPHY_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23718_ _23753_/CLK _20523_/Y HRESETn VGND VGND VPWR VPWR _20520_/A sky130_fd_sc_hd__dfrtp_4
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24698_ _24698_/CLK _24698_/D HRESETn VGND VGND VPWR VPWR _24698_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24969__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14451_ _21657_/A VGND VGND VPWR VPWR _14524_/B sky130_fd_sc_hd__buf_2
XPHY_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11663_ _11663_/A VGND VGND VPWR VPWR _11663_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23649_ _24823_/CLK _23649_/D HRESETn VGND VGND VPWR VPWR _23649_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13402_/A VGND VGND VPWR VPWR _21700_/A sky130_fd_sc_hd__inv_2
XANTENNA__22275__B _21300_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17170_ _17186_/A VGND VGND VPWR VPWR _17170_/Y sky130_fd_sc_hd__inv_2
XPHY_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14382_ _13438_/Y _14382_/B VGND VGND VPWR VPWR _14383_/B sky130_fd_sc_hd__or2_4
XPHY_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11594_ _16096_/A VGND VGND VPWR VPWR _11594_/X sky130_fd_sc_hd__buf_2
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16121_ _16121_/A VGND VGND VPWR VPWR _16121_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_114_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_229_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13333_ _13333_/A VGND VGND VPWR VPWR _20818_/A sky130_fd_sc_hd__buf_2
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24551__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16052_ _16071_/A VGND VGND VPWR VPWR _16052_/X sky130_fd_sc_hd__buf_2
X_13264_ _13232_/A _13260_/X _13264_/C VGND VGND VPWR VPWR _13264_/X sky130_fd_sc_hd__or3_4
XFILLER_68_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15003_ _15003_/A _15003_/B _15123_/B VGND VGND VPWR VPWR _15012_/A sky130_fd_sc_hd__or3_4
X_12215_ _12215_/A VGND VGND VPWR VPWR _12215_/Y sky130_fd_sc_hd__inv_2
X_13195_ _13120_/X _18863_/A VGND VGND VPWR VPWR _13195_/X sky130_fd_sc_hd__or2_4
XFILLER_9_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19811_ _19801_/A _18067_/A _11643_/A _23199_/Q _19802_/A VGND VGND VPWR VPWR _19811_/X
+ sky130_fd_sc_hd__a32o_4
X_12146_ _24565_/Q VGND VGND VPWR VPWR _12146_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22719__A2 _22536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19742_ _19742_/A VGND VGND VPWR VPWR _21824_/B sky130_fd_sc_hd__inv_2
XANTENNA__19045__B1 _18953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12077_ _25108_/Q _12075_/Y _12185_/A _12089_/A VGND VGND VPWR VPWR _12077_/X sky130_fd_sc_hd__a2bb2o_4
X_16954_ _16921_/D VGND VGND VPWR VPWR _16954_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12322__A _12322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15905_ _15904_/Y _15900_/X _15801_/X _15900_/X VGND VGND VPWR VPWR _15905_/X sky130_fd_sc_hd__a2bb2o_4
X_19673_ _19680_/A VGND VGND VPWR VPWR _19673_/X sky130_fd_sc_hd__buf_2
X_16885_ _16885_/A _16885_/B VGND VGND VPWR VPWR _16885_/X sky130_fd_sc_hd__or2_4
XANTENNA__15606__B1 _11563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18624_ _18624_/A VGND VGND VPWR VPWR _18624_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_52_0_HCLK clkbuf_8_53_0_HCLK/A VGND VGND VPWR VPWR _23085_/CLK sky130_fd_sc_hd__clkbuf_1
X_15836_ _24423_/Q VGND VGND VPWR VPWR _15836_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20896__D _20896_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18555_ _18552_/A _18552_/B VGND VGND VPWR VPWR _18555_/Y sky130_fd_sc_hd__nand2_4
XFILLER_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12979_ _12863_/Y _12974_/B VGND VGND VPWR VPWR _12992_/B sky130_fd_sc_hd__or2_4
X_15767_ _15750_/Y VGND VGND VPWR VPWR _15767_/X sky130_fd_sc_hd__buf_2
XFILLER_18_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17359__B1 _17336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22352__B1 _22351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18944__A _18943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17506_ _17505_/X VGND VGND VPWR VPWR _17508_/B sky130_fd_sc_hd__inv_2
XANTENNA__19657__A1_N _19656_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14718_ _15085_/A _24093_/Q _15085_/A _24093_/Q VGND VGND VPWR VPWR _14718_/X sky130_fd_sc_hd__a2bb2o_4
X_18486_ _18430_/Y _18486_/B _18507_/B VGND VGND VPWR VPWR _18495_/D sky130_fd_sc_hd__or3_4
X_15698_ _15695_/A VGND VGND VPWR VPWR _15698_/X sky130_fd_sc_hd__buf_2
XFILLER_61_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17437_ _17320_/A _17435_/X VGND VGND VPWR VPWR _17438_/B sky130_fd_sc_hd__or2_4
XFILLER_53_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14649_ _14636_/X _14648_/Y _24727_/Q _14636_/X VGND VGND VPWR VPWR _14649_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12992__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24639__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22655__A1 _23961_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17368_ _17622_/B _17363_/Y _17368_/C VGND VGND VPWR VPWR _17368_/X sky130_fd_sc_hd__or3_4
XFILLER_119_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19107_ _19105_/Y _19101_/X _19041_/X _19106_/X VGND VGND VPWR VPWR _19107_/X sky130_fd_sc_hd__a2bb2o_4
X_16319_ _16318_/Y _16314_/X _16246_/X _16314_/X VGND VGND VPWR VPWR _24249_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17299_ _17510_/B VGND VGND VPWR VPWR _17505_/C sky130_fd_sc_hd__buf_2
XANTENNA__24292__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22913__B _22015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19038_ _18739_/X VGND VGND VPWR VPWR _19038_/X sky130_fd_sc_hd__buf_2
XANTENNA__15688__A3 _15499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24221__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14896__B2 _24271_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_19_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_115_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21000_ _21007_/A _21000_/B _20999_/X VGND VGND VPWR VPWR _21000_/X sky130_fd_sc_hd__and3_4
XFILLER_138_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15527__B _15531_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15845__B1 _11548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19036__B1 _18901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22951_ _22730_/A _22951_/B VGND VGND VPWR VPWR _22951_/Y sky130_fd_sc_hd__nor2_4
XFILLER_110_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21902_ _20239_/A _14016_/X _14081_/A _20802_/X VGND VGND VPWR VPWR _21905_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25080__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22882_ _24249_/Q _21553_/X _20780_/X _22881_/X VGND VGND VPWR VPWR _22882_/X sky130_fd_sc_hd__a211o_4
X_24621_ _24587_/CLK _15305_/X HRESETn VGND VGND VPWR VPWR _11951_/B sky130_fd_sc_hd__dfrtp_4
X_21833_ _20978_/A _19559_/Y _17642_/Y VGND VGND VPWR VPWR _21833_/X sky130_fd_sc_hd__o21a_4
XFILLER_43_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24552_ _24566_/CLK _15516_/X HRESETn VGND VGND VPWR VPWR _24552_/Q sky130_fd_sc_hd__dfrtp_4
X_21764_ _21764_/A _21761_/X _21763_/X VGND VGND VPWR VPWR _21764_/X sky130_fd_sc_hd__and3_4
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22376__A _22376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23503_ _23511_/CLK _18965_/X VGND VGND VPWR VPWR _18963_/A sky130_fd_sc_hd__dfxtp_4
X_20715_ _20715_/A _20713_/Y VGND VGND VPWR VPWR _20715_/Y sky130_fd_sc_hd__nor2_4
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24483_ _24483_/CLK _24483_/D HRESETn VGND VGND VPWR VPWR _24483_/Q sky130_fd_sc_hd__dfrtp_4
X_21695_ _13468_/A _19279_/Y _21696_/A _21251_/A VGND VGND VPWR VPWR _21695_/X sky130_fd_sc_hd__o22a_4
XFILLER_106_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23434_ _25067_/CLK _19158_/X VGND VGND VPWR VPWR _23434_/Q sky130_fd_sc_hd__dfxtp_4
X_20646_ _20621_/X _20645_/Y _16505_/A _20624_/X VGND VGND VPWR VPWR _23747_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24309__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23365_ _23374_/CLK _23365_/D VGND VGND VPWR VPWR _23365_/Q sky130_fd_sc_hd__dfxtp_4
X_20577_ _21729_/A _20574_/X _20562_/X _20576_/X VGND VGND VPWR VPWR _20578_/A sky130_fd_sc_hd__o22a_4
XFILLER_20_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12407__A _12406_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25104_ _25112_/CLK _12297_/X HRESETn VGND VGND VPWR VPWR _12113_/A sky130_fd_sc_hd__dfrtp_4
X_22316_ _22225_/X _22313_/X _22231_/X _22315_/X VGND VGND VPWR VPWR _22317_/B sky130_fd_sc_hd__o22a_4
X_23296_ _23385_/CLK _19549_/X VGND VGND VPWR VPWR _23296_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20624__A _20651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12843__A2_N _22463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22949__A2 _21896_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25035_ _24435_/CLK _12898_/Y HRESETn VGND VGND VPWR VPWR _22980_/A sky130_fd_sc_hd__dfrtp_4
X_22247_ _23025_/B _22246_/X _22197_/X _24405_/Q _20866_/X VGND VGND VPWR VPWR _22248_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_69_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19275__B1 _19227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12000_ _11999_/Y _11995_/X _11620_/X _11995_/X VGND VGND VPWR VPWR _25143_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11965__B _11956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22178_ _22178_/A VGND VGND VPWR VPWR _22178_/X sky130_fd_sc_hd__buf_2
X_21129_ _17631_/Y VGND VGND VPWR VPWR _21339_/A sky130_fd_sc_hd__buf_2
XANTENNA__17933__A _17716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23944__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25168__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13951_ _13950_/X VGND VGND VPWR VPWR _13952_/A sky130_fd_sc_hd__buf_2
XANTENNA__16549__A _16530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11981__A _13398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12902_ _12812_/Y _12899_/X VGND VGND VPWR VPWR _12902_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_39_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_79_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13882_ _20271_/A _20164_/A _13887_/A _13898_/A VGND VGND VPWR VPWR _13885_/A sky130_fd_sc_hd__o22a_4
X_16670_ _16652_/X _16653_/X _15706_/X _24096_/Q _16647_/X VGND VGND VPWR VPWR _16670_/X
+ sky130_fd_sc_hd__a32o_4
X_12833_ _12880_/B VGND VGND VPWR VPWR _12833_/X sky130_fd_sc_hd__buf_2
X_15621_ _15604_/A VGND VGND VPWR VPWR _15621_/X sky130_fd_sc_hd__buf_2
X_24819_ _24788_/CLK _14214_/X HRESETn VGND VGND VPWR VPWR _14211_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18764__A _18763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18340_ _23844_/Q VGND VGND VPWR VPWR _18442_/A sky130_fd_sc_hd__buf_2
X_12764_ _12629_/X _12765_/B VGND VGND VPWR VPWR _12766_/A sky130_fd_sc_hd__nand2_4
X_15552_ _19828_/A VGND VGND VPWR VPWR _19455_/A sky130_fd_sc_hd__buf_2
XANTENNA__22885__A1 _21561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _11698_/D _11714_/X _11703_/X VGND VGND VPWR VPWR _11715_/X sky130_fd_sc_hd__o21a_4
X_14503_ _14502_/Y _14480_/A _21751_/A _14484_/X VGND VGND VPWR VPWR _14517_/B sky130_fd_sc_hd__o22a_4
XFILLER_76_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _15460_/X VGND VGND VPWR VPWR _15483_/X sky130_fd_sc_hd__buf_2
X_18271_ _18270_/X VGND VGND VPWR VPWR _18271_/Y sky130_fd_sc_hd__inv_2
X_12695_ _12654_/X _12663_/B _12612_/Y VGND VGND VPWR VPWR _12695_/X sky130_fd_sc_hd__o21a_4
XPHY_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24732__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _17197_/B _17222_/B VGND VGND VPWR VPWR _17222_/Y sky130_fd_sc_hd__nor2_4
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11646_ _11645_/X VGND VGND VPWR VPWR _11708_/B sky130_fd_sc_hd__inv_2
X_14434_ _14434_/A _14433_/X VGND VGND VPWR VPWR _14435_/D sky130_fd_sc_hd__and2_4
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14365_ HSEL VGND VGND VPWR VPWR _14366_/A sky130_fd_sc_hd__buf_2
X_17153_ _17129_/A _17153_/B _17152_/Y VGND VGND VPWR VPWR _24033_/D sky130_fd_sc_hd__and3_4
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11577_ _11541_/X VGND VGND VPWR VPWR _11577_/X sky130_fd_sc_hd__buf_2
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17513__B1 _16748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13316_ _13316_/A _23319_/Q VGND VGND VPWR VPWR _13317_/C sky130_fd_sc_hd__or2_4
X_16104_ _24333_/Q VGND VGND VPWR VPWR _22232_/A sky130_fd_sc_hd__inv_2
X_17084_ _17026_/B _17077_/X _17083_/X _17079_/Y VGND VGND VPWR VPWR _17085_/A sky130_fd_sc_hd__a211o_4
X_14296_ _14295_/Y _14293_/X _14209_/X _14293_/X VGND VGND VPWR VPWR _14296_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13247_ _13247_/A _13243_/X _13246_/X VGND VGND VPWR VPWR _13247_/X sky130_fd_sc_hd__or3_4
X_16035_ _16035_/A _16035_/B _16027_/X _16034_/X VGND VGND VPWR VPWR _16035_/X sky130_fd_sc_hd__or4_4
XANTENNA__15628__A _15604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13178_ _13316_/A _13178_/B VGND VGND VPWR VPWR _13178_/X sky130_fd_sc_hd__or2_4
XFILLER_123_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11561__B1 _25211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12129_ _12129_/A VGND VGND VPWR VPWR _12237_/A sky130_fd_sc_hd__inv_2
XFILLER_96_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17986_ _17982_/X _15430_/X _16096_/A _23922_/Q _17983_/X VGND VGND VPWR VPWR _23922_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_112_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12105__A2 _24552_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19725_ _21459_/B _19718_/X _19724_/X _19718_/X VGND VGND VPWR VPWR _19725_/X sky130_fd_sc_hd__a2bb2o_4
X_16937_ _16771_/Y _16937_/B VGND VGND VPWR VPWR _16937_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12368__A1_N _12498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19656_ _19656_/A VGND VGND VPWR VPWR _19656_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11864__A1 _21188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16868_ _16879_/A _16841_/X _16819_/Y VGND VGND VPWR VPWR _16868_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16252__B1 _16251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18607_ _18607_/A VGND VGND VPWR VPWR _18607_/X sky130_fd_sc_hd__buf_2
X_15819_ _11529_/A VGND VGND VPWR VPWR _22933_/B sky130_fd_sc_hd__buf_2
XFILLER_52_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19587_ _19587_/A VGND VGND VPWR VPWR _21383_/B sky130_fd_sc_hd__inv_2
X_16799_ _15899_/Y _16835_/A _24423_/Q _16853_/A VGND VGND VPWR VPWR _16804_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14802__B2 _14801_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18538_ _18532_/A _18536_/X _18537_/Y VGND VGND VPWR VPWR _23822_/D sky130_fd_sc_hd__o21a_4
XFILLER_94_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19741__B2 _19738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18469_ _18469_/A _18468_/X VGND VGND VPWR VPWR _18470_/B sky130_fd_sc_hd__or2_4
XANTENNA__24473__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20500_ _20498_/Y _20495_/X _20499_/X VGND VGND VPWR VPWR _20500_/X sky130_fd_sc_hd__o21a_4
XFILLER_18_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21480_ _21476_/X _21479_/X _21930_/A VGND VGND VPWR VPWR _21480_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12306__A1_N _12305_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22924__A _14777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24402__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20431_ _15398_/Y _20416_/X _20425_/X _20430_/X VGND VGND VPWR VPWR _20431_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23150_ _23596_/CLK _23150_/D VGND VGND VPWR VPWR _23150_/Q sky130_fd_sc_hd__dfxtp_4
X_20362_ _20361_/X VGND VGND VPWR VPWR _23670_/D sky130_fd_sc_hd__inv_2
XANTENNA__14947__A2_N _24278_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22101_ _20962_/A _22101_/B _22100_/X VGND VGND VPWR VPWR _22101_/X sky130_fd_sc_hd__and3_4
X_23081_ _23908_/CLK _20125_/X VGND VGND VPWR VPWR _23081_/Q sky130_fd_sc_hd__dfxtp_4
X_20293_ _20293_/A _20292_/Y _20278_/X VGND VGND VPWR VPWR _20293_/X sky130_fd_sc_hd__and3_4
XANTENNA__15530__A2 _15319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22032_ _22006_/B _22030_/X _21881_/A _22031_/X VGND VGND VPWR VPWR _22032_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20811__B1 _20801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17753__A _17918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16491__B1 _16153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18175__A1_N _16080_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21275__A _21275_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23983_ _23990_/CLK _23983_/D HRESETn VGND VGND VPWR VPWR _17430_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21706__C _21653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16369__A _16369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21693__A1_N _15430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22934_ _15331_/Y _22870_/B VGND VGND VPWR VPWR _22934_/X sky130_fd_sc_hd__and2_4
XFILLER_84_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22865_ _24350_/Q _22311_/A _22864_/X VGND VGND VPWR VPWR _22865_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15597__A2 _15582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17991__B1 _22215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21816_ _20966_/A _19672_/Y VGND VGND VPWR VPWR _21816_/X sky130_fd_sc_hd__or2_4
X_24604_ _24604_/CLK _15354_/X HRESETn VGND VGND VPWR VPWR _15352_/A sky130_fd_sc_hd__dfrtp_4
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22796_ _12101_/Y _21042_/A _12332_/Y _22238_/X VGND VGND VPWR VPWR _22796_/X sky130_fd_sc_hd__o22a_4
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19732__B2 _19727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24535_ _25061_/CLK _15564_/X HRESETn VGND VGND VPWR VPWR _19835_/A sky130_fd_sc_hd__dfrtp_4
X_21747_ _19265_/Y _21082_/B _21582_/X _21746_/X VGND VGND VPWR VPWR _21747_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15816__A1_N _15712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11500_ _11938_/A _14013_/B VGND VGND VPWR VPWR _11500_/X sky130_fd_sc_hd__or2_4
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12480_ _12460_/A _12480_/B _12479_/Y VGND VGND VPWR VPWR _25088_/D sky130_fd_sc_hd__and3_4
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24466_ _23442_/CLK _24466_/D HRESETn VGND VGND VPWR VPWR _24466_/Q sky130_fd_sc_hd__dfrtp_4
X_21678_ _21202_/A _21678_/B _21678_/C VGND VGND VPWR VPWR _21678_/X sky130_fd_sc_hd__and3_4
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22834__A _24315_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24143__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23417_ _23416_/CLK _19205_/X VGND VGND VPWR VPWR _23417_/Q sky130_fd_sc_hd__dfxtp_4
X_20629_ _20621_/X _20628_/Y _24174_/Q _20624_/X VGND VGND VPWR VPWR _23743_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24397_ _24587_/CLK _15905_/X HRESETn VGND VGND VPWR VPWR _24397_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14150_ _14149_/X VGND VGND VPWR VPWR _14150_/X sky130_fd_sc_hd__buf_2
XANTENNA__12583__A2 _12582_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23348_ _23350_/CLK _23348_/D VGND VGND VPWR VPWR _13146_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_138_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13101_ _13247_/A _13095_/X _13100_/X VGND VGND VPWR VPWR _13101_/X sky130_fd_sc_hd__or3_4
XFILLER_3_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14081_ _14081_/A VGND VGND VPWR VPWR _14081_/Y sky130_fd_sc_hd__inv_2
X_23279_ _23303_/CLK _19593_/X VGND VGND VPWR VPWR _19592_/A sky130_fd_sc_hd__dfxtp_4
X_13032_ _18085_/A _13032_/B VGND VGND VPWR VPWR _13032_/X sky130_fd_sc_hd__or2_4
X_25018_ _24523_/CLK _25018_/D HRESETn VGND VGND VPWR VPWR _22396_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__11695__B _11694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11543__B1 _11540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17840_ _17968_/A _17840_/B _17839_/X VGND VGND VPWR VPWR _17840_/X sky130_fd_sc_hd__and3_4
XFILLER_43_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16482__B1 _16141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17771_ _17729_/A VGND VGND VPWR VPWR _17878_/A sky130_fd_sc_hd__buf_2
XANTENNA__17382__B _17270_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14983_ _14882_/A _14881_/X _14990_/A _14982_/X VGND VGND VPWR VPWR _14983_/X sky130_fd_sc_hd__or4_4
XANTENNA__12099__B2 _12098_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16279__A HWDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19510_ _19509_/X VGND VGND VPWR VPWR _19510_/Y sky130_fd_sc_hd__inv_2
X_16722_ _23947_/Q VGND VGND VPWR VPWR _21839_/A sky130_fd_sc_hd__inv_2
X_13934_ _13934_/A _13934_/B _13934_/C VGND VGND VPWR VPWR _13935_/A sky130_fd_sc_hd__or3_4
XFILLER_74_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24984__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19441_ _19440_/Y VGND VGND VPWR VPWR _19441_/X sky130_fd_sc_hd__buf_2
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20030__B2 _20027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16653_ _16625_/A VGND VGND VPWR VPWR _16653_/X sky130_fd_sc_hd__buf_2
X_13865_ _13864_/X VGND VGND VPWR VPWR _13865_/Y sky130_fd_sc_hd__inv_2
X_15604_ _15604_/A VGND VGND VPWR VPWR _15604_/X sky130_fd_sc_hd__buf_2
X_12816_ _22187_/A VGND VGND VPWR VPWR _12816_/Y sky130_fd_sc_hd__inv_2
X_19372_ _19372_/A VGND VGND VPWR VPWR _19372_/Y sky130_fd_sc_hd__inv_2
X_16584_ _16584_/A VGND VGND VPWR VPWR _16584_/X sky130_fd_sc_hd__buf_2
XFILLER_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13796_ _13796_/A _13735_/A VGND VGND VPWR VPWR _13797_/C sky130_fd_sc_hd__and2_4
XFILLER_128_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_126_0_HCLK clkbuf_7_63_0_HCLK/X VGND VGND VPWR VPWR _23859_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18323_ _18302_/X _18323_/B _18319_/X VGND VGND VPWR VPWR _23850_/D sky130_fd_sc_hd__and3_4
X_15535_ _14369_/B _14435_/D _15438_/A _14431_/A VGND VGND VPWR VPWR _15535_/X sky130_fd_sc_hd__and4_4
X_12747_ _12749_/A _12747_/B _12746_/Y VGND VGND VPWR VPWR _12747_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_189_0_HCLK clkbuf_7_94_0_HCLK/X VGND VGND VPWR VPWR _24488_/CLK sky130_fd_sc_hd__clkbuf_1
X_18254_ _18226_/A _18250_/X _18253_/Y VGND VGND VPWR VPWR _23869_/D sky130_fd_sc_hd__and3_4
X_12678_ _12605_/Y _12677_/X VGND VGND VPWR VPWR _12694_/B sky130_fd_sc_hd__or2_4
X_15466_ _15466_/A VGND VGND VPWR VPWR _15466_/X sky130_fd_sc_hd__buf_2
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17205_ _16376_/A VGND VGND VPWR VPWR _17205_/X sky130_fd_sc_hd__buf_2
X_11629_ HWDATA[3] VGND VGND VPWR VPWR _11630_/A sky130_fd_sc_hd__buf_2
X_14417_ _14377_/A _14377_/B VGND VGND VPWR VPWR _14417_/X sky130_fd_sc_hd__or2_4
XFILLER_30_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18185_ _18178_/X _18180_/X _18182_/X _18185_/D VGND VGND VPWR VPWR _18191_/C sky130_fd_sc_hd__or4_4
X_15397_ _15395_/Y _15396_/X _15279_/X _15396_/X VGND VGND VPWR VPWR _15397_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15760__A2 _15740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17136_ _17135_/X VGND VGND VPWR VPWR _17137_/B sky130_fd_sc_hd__inv_2
X_14348_ _20271_/A _13899_/B VGND VGND VPWR VPWR _14348_/X sky130_fd_sc_hd__and2_4
XANTENNA__15358__A _15401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23866__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14279_ _24794_/Q VGND VGND VPWR VPWR _14279_/Y sky130_fd_sc_hd__inv_2
X_17067_ _17067_/A _17046_/X VGND VGND VPWR VPWR _17070_/B sky130_fd_sc_hd__or2_4
XFILLER_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14262__A _24801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16018_ _16014_/A _16016_/X _16012_/X _16017_/Y VGND VGND VPWR VPWR _24358_/D sky130_fd_sc_hd__o22a_4
XFILLER_131_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25019__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22794__B1 _21882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21807__B _21807_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17969_ _17969_/A _17969_/B _17968_/X VGND VGND VPWR VPWR _17970_/C sky130_fd_sc_hd__or3_4
XFILLER_61_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19708_ _19530_/X _18025_/D _19236_/X VGND VGND VPWR VPWR _19709_/A sky130_fd_sc_hd__or3_4
X_20980_ _20980_/A _20978_/X _20980_/C VGND VGND VPWR VPWR _20980_/X sky130_fd_sc_hd__and3_4
XANTENNA__12510__A _12408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19639_ _21145_/B _19636_/X _19617_/X _19636_/X VGND VGND VPWR VPWR _23264_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_22_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16917__A _16936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24654__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_85_0_HCLK clkbuf_6_42_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_85_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__22849__A1 _23020_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22650_ _21050_/Y VGND VGND VPWR VPWR _22651_/B sky130_fd_sc_hd__buf_2
XANTENNA__22849__B2 _20833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21601_ _21600_/X VGND VGND VPWR VPWR _21601_/Y sky130_fd_sc_hd__inv_2
X_22581_ _22351_/A VGND VGND VPWR VPWR _22581_/X sky130_fd_sc_hd__buf_2
XFILLER_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24320_ _24289_/CLK _24320_/D HRESETn VGND VGND VPWR VPWR _22999_/A sky130_fd_sc_hd__dfrtp_4
X_21532_ _20892_/X _21531_/X _24944_/Q _22548_/A VGND VGND VPWR VPWR _21532_/X sky130_fd_sc_hd__o22a_4
XFILLER_138_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24251_ _24192_/CLK _16315_/X HRESETn VGND VGND VPWR VPWR _16312_/A sky130_fd_sc_hd__dfrtp_4
X_21463_ _21333_/A _21463_/B VGND VGND VPWR VPWR _21463_/X sky130_fd_sc_hd__or2_4
XANTENNA__16652__A _16624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21445__A2_N _11503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14886__A2_N _24286_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22373__B _22524_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23202_ _23990_/CLK _23202_/D VGND VGND VPWR VPWR _13205_/B sky130_fd_sc_hd__dfxtp_4
X_20414_ _20414_/A _13516_/X VGND VGND VPWR VPWR _20414_/X sky130_fd_sc_hd__or2_4
X_24182_ _24182_/CLK _16496_/X HRESETn VGND VGND VPWR VPWR _16495_/A sky130_fd_sc_hd__dfrtp_4
X_21394_ _21394_/A _21394_/B _21394_/C VGND VGND VPWR VPWR _21394_/X sky130_fd_sc_hd__and3_4
XFILLER_49_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23133_ _23133_/CLK _19994_/X VGND VGND VPWR VPWR _23133_/Q sky130_fd_sc_hd__dfxtp_4
X_20345_ _20345_/A _17187_/X VGND VGND VPWR VPWR _20345_/X sky130_fd_sc_hd__and2_4
XANTENNA__19963__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21037__B1 _24546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23064_ _23624_/CLK scl_oen_o_S4 VGND VGND VPWR VPWR _20702_/A sky130_fd_sc_hd__dfxtp_4
X_20276_ _20276_/A VGND VGND VPWR VPWR _20276_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20902__A _11720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22015_ _20786_/A VGND VGND VPWR VPWR _22015_/X sky130_fd_sc_hd__buf_2
XFILLER_66_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15267__A1 _14100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14900__A _14900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11980_ _11980_/A VGND VGND VPWR VPWR _11980_/Y sky130_fd_sc_hd__inv_2
X_23966_ _24378_/CLK _23966_/D HRESETn VGND VGND VPWR VPWR _22782_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21745__D1 _21744_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22917_ _16621_/A _22916_/X _22839_/X _24573_/Q _21694_/X VGND VGND VPWR VPWR _22917_/X
+ sky130_fd_sc_hd__a32o_4
X_23897_ _23979_/CLK _18071_/Y HRESETn VGND VGND VPWR VPWR _23897_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24395__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13650_ _22483_/A _13649_/X _11581_/X _13649_/X VGND VGND VPWR VPWR _24940_/D sky130_fd_sc_hd__a2bb2o_4
X_22848_ _24493_/Q _13618_/A VGND VGND VPWR VPWR _22848_/X sky130_fd_sc_hd__or2_4
XANTENNA__24324__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _12644_/D _24516_/Q _12644_/D _24516_/Q VGND VGND VPWR VPWR _12601_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22304__A3 _22251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13581_ _13564_/A _13563_/X VGND VGND VPWR VPWR _13581_/Y sky130_fd_sc_hd__nand2_4
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22779_ _22779_/A _22147_/A VGND VGND VPWR VPWR _22779_/X sky130_fd_sc_hd__and2_4
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12532_ _12389_/X _12535_/B _12427_/X VGND VGND VPWR VPWR _12532_/Y sky130_fd_sc_hd__a21oi_4
X_15320_ HWDATA[31] VGND VGND VPWR VPWR _15320_/X sky130_fd_sc_hd__buf_2
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24518_ _24483_/CLK _24518_/D HRESETn VGND VGND VPWR VPWR _24518_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12463_ _12463_/A VGND VGND VPWR VPWR _12463_/Y sky130_fd_sc_hd__inv_2
X_15251_ _15251_/A _15251_/B VGND VGND VPWR VPWR _15251_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__19469__B1 _17993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24449_ _24432_/CLK _24449_/D HRESETn VGND VGND VPWR VPWR _24449_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16562__A _21590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15742__A2 _15740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14202_ _14201_/X VGND VGND VPWR VPWR _14202_/X sky130_fd_sc_hd__buf_2
X_15182_ _24665_/Q _15182_/B VGND VGND VPWR VPWR _15183_/C sky130_fd_sc_hd__or2_4
XANTENNA__20039__A2_N _20036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12394_ _25076_/Q VGND VGND VPWR VPWR _12408_/C sky130_fd_sc_hd__inv_2
XFILLER_138_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14133_ _24846_/Q _14122_/X _24845_/Q _14127_/X VGND VGND VPWR VPWR _14133_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23017__A1 _24286_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19990_ _19989_/X VGND VGND VPWR VPWR _19990_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25183__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14064_ _14064_/A VGND VGND VPWR VPWR _14064_/Y sky130_fd_sc_hd__inv_2
X_18941_ _18940_/Y _18935_/X _18828_/X _18935_/A VGND VGND VPWR VPWR _18941_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21908__A _17629_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20812__A _22564_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25112__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22776__B1 _14729_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13015_ _13078_/A VGND VGND VPWR VPWR _13016_/A sky130_fd_sc_hd__buf_2
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18872_ _17681_/B VGND VGND VPWR VPWR _18872_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15906__A _24396_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15258__A1 _14100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17823_ _17738_/A _17823_/B _17822_/X VGND VGND VPWR VPWR _17824_/C sky130_fd_sc_hd__or3_4
XFILLER_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16960__A2_N _24058_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22528__B1 _17041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17754_ _17742_/A VGND VGND VPWR VPWR _17927_/A sky130_fd_sc_hd__buf_2
XFILLER_94_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14966_ _24680_/Q VGND VGND VPWR VPWR _14966_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14481__A2 _14475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16705_ _17490_/B VGND VGND VPWR VPWR _17595_/C sky130_fd_sc_hd__buf_2
X_13917_ _13916_/X _14361_/B _13896_/X _24898_/Q _13911_/X VGND VGND VPWR VPWR _13917_/X
+ sky130_fd_sc_hd__a32o_4
X_17685_ _17698_/A _17685_/B VGND VGND VPWR VPWR _17685_/X sky130_fd_sc_hd__or2_4
XFILLER_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14897_ _14897_/A VGND VGND VPWR VPWR _14897_/Y sky130_fd_sc_hd__inv_2
X_19424_ HWDATA[5] VGND VGND VPWR VPWR _19424_/X sky130_fd_sc_hd__buf_2
XANTENNA__15641__A _22218_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22458__B _22238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16636_ _14729_/Y _16632_/X HWDATA[24] _16632_/X VGND VGND VPWR VPWR _16636_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14769__B1 _14712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13848_ _13812_/X _13843_/Y _13844_/Y _13813_/Y _13847_/Y VGND VGND VPWR VPWR _13848_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24065__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19355_ _19349_/Y VGND VGND VPWR VPWR _19355_/X sky130_fd_sc_hd__buf_2
XFILLER_62_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16567_ _15799_/X _16276_/X _15743_/X _24156_/Q _16566_/X VGND VGND VPWR VPWR _16567_/X
+ sky130_fd_sc_hd__a32o_4
X_13779_ _13764_/X _13770_/B _13716_/D _13779_/D VGND VGND VPWR VPWR _13779_/X sky130_fd_sc_hd__and4_4
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18306_ _18312_/A _18312_/B VGND VGND VPWR VPWR _18307_/B sky130_fd_sc_hd__or2_4
X_15518_ _15470_/Y VGND VGND VPWR VPWR _15518_/X sky130_fd_sc_hd__buf_2
X_19286_ _23389_/Q VGND VGND VPWR VPWR _21928_/B sky130_fd_sc_hd__inv_2
X_16498_ _16479_/A VGND VGND VPWR VPWR _16499_/A sky130_fd_sc_hd__buf_2
X_18237_ _18559_/B VGND VGND VPWR VPWR _18237_/X sky130_fd_sc_hd__buf_2
XFILLER_50_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15449_ _15449_/A _15449_/B VGND VGND VPWR VPWR _15453_/A sky130_fd_sc_hd__and2_4
XFILLER_129_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19287__A2_N _19284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21267__B1 _25192_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18168_ _18322_/A VGND VGND VPWR VPWR _18216_/A sky130_fd_sc_hd__inv_2
XFILLER_11_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17119_ _17040_/A _17116_/X VGND VGND VPWR VPWR _17120_/C sky130_fd_sc_hd__or2_4
XFILLER_89_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16289__A3 _15706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18099_ _18099_/A VGND VGND VPWR VPWR _18099_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20130_ _13923_/B _13923_/C VGND VGND VPWR VPWR _20131_/A sky130_fd_sc_hd__or2_4
XANTENNA__21818__A _20972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22767__B1 _15849_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20061_ _20058_/Y _20060_/X _19424_/X _20060_/X VGND VGND VPWR VPWR _20061_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22519__B1 _24518_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16997__B2 _24039_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13336__A _13335_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24835__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23820_ _23826_/CLK _18542_/X HRESETn VGND VGND VPWR VPWR _23820_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21553__A _21553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23751_ _24112_/CLK _20662_/X HRESETn VGND VGND VPWR VPWR _23751_/Q sky130_fd_sc_hd__dfrtp_4
X_20963_ _21130_/A VGND VGND VPWR VPWR _20967_/A sky130_fd_sc_hd__buf_2
XFILLER_22_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16647__A _16627_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21742__B2 _21400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22702_ _22702_/A _22702_/B VGND VGND VPWR VPWR _22702_/X sky130_fd_sc_hd__and2_4
X_23682_ _24769_/CLK _23681_/Q HRESETn VGND VGND VPWR VPWR _23682_/Q sky130_fd_sc_hd__dfrtp_4
X_20894_ _22311_/A _20884_/X _20890_/X _20891_/X _20893_/X VGND VGND VPWR VPWR _20894_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_13_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22633_ _22633_/A _22703_/B VGND VGND VPWR VPWR _22633_/X sky130_fd_sc_hd__or2_4
XFILLER_80_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22564_ _22564_/A _22564_/B VGND VGND VPWR VPWR _22564_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_172_0_HCLK clkbuf_7_86_0_HCLK/X VGND VGND VPWR VPWR _23135_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18371__B1 _16400_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21515_ _21224_/A _21513_/X _21515_/C VGND VGND VPWR VPWR _21515_/X sky130_fd_sc_hd__and3_4
XANTENNA__23788__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24303_ _24037_/CLK _24303_/D HRESETn VGND VGND VPWR VPWR _16183_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17478__A _22979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22495_ _22495_/A _22486_/Y _22490_/Y _22495_/D VGND VGND VPWR VPWR _22495_/X sky130_fd_sc_hd__or4_4
Xclkbuf_8_29_0_HCLK clkbuf_8_29_0_HCLK/A VGND VGND VPWR VPWR _24928_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_6_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21258__B1 _21256_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23717__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24234_ _24201_/CLK _16357_/X HRESETn VGND VGND VPWR VPWR _24234_/Q sky130_fd_sc_hd__dfrtp_4
X_21446_ _24795_/Q _20931_/X _21443_/X _21444_/X _21445_/X VGND VGND VPWR VPWR _21446_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_119_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24165_ _24167_/CLK _16538_/X HRESETn VGND VGND VPWR VPWR _16537_/A sky130_fd_sc_hd__dfrtp_4
X_21377_ _21214_/A _21377_/B VGND VGND VPWR VPWR _21377_/X sky130_fd_sc_hd__or2_4
XANTENNA__12415__A _12415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23116_ _23293_/CLK _23116_/D VGND VGND VPWR VPWR _20038_/A sky130_fd_sc_hd__dfxtp_4
X_20328_ _20328_/A VGND VGND VPWR VPWR _20328_/Y sky130_fd_sc_hd__inv_2
X_24096_ _24094_/CLK _16670_/X HRESETn VGND VGND VPWR VPWR _24096_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22758__B1 _24568_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23047_ VGND VGND VPWR VPWR _23047_/HI IRQ[15] sky130_fd_sc_hd__conb_1
X_20259_ _23766_/Q _20265_/B _20247_/X VGND VGND VPWR VPWR _20259_/X sky130_fd_sc_hd__a21o_4
XFILLER_77_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16437__B1 _16087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24576__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14820_ _14813_/X _14820_/B _14817_/X _14819_/X VGND VGND VPWR VPWR _14820_/X sky130_fd_sc_hd__or4_4
XFILLER_44_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22559__A _15653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24998_ _24998_/CLK _13257_/X HRESETn VGND VGND VPWR VPWR _24998_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24505__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21463__A _21333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14751_ _14751_/A VGND VGND VPWR VPWR _14751_/Y sky130_fd_sc_hd__inv_2
X_11963_ _22564_/B VGND VGND VPWR VPWR _11964_/A sky130_fd_sc_hd__buf_2
XFILLER_56_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23949_ _23949_/CLK _23949_/D HRESETn VGND VGND VPWR VPWR _16704_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20536__A2 _20416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14778__A2_N _24097_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22930__B1 _22858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22278__B _22188_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13702_ _24917_/Q _13686_/X _24916_/Q _13681_/X VGND VGND VPWR VPWR _13702_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15461__A _15460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17470_ _17454_/X _17458_/Y VGND VGND VPWR VPWR _17470_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__21182__B _20827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11894_ _11894_/A VGND VGND VPWR VPWR _11894_/Y sky130_fd_sc_hd__inv_2
X_14682_ _14682_/A VGND VGND VPWR VPWR _14682_/X sky130_fd_sc_hd__buf_2
XFILLER_72_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16421_ _16426_/A VGND VGND VPWR VPWR _16421_/X sky130_fd_sc_hd__buf_2
X_13633_ _13622_/Y _13631_/X _13632_/X _13631_/X VGND VGND VPWR VPWR _13633_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22289__A2 _22230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19140_ _19139_/Y _19137_/X _19095_/X _19137_/X VGND VGND VPWR VPWR _19140_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14701__A2_N _14699_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16352_ _16364_/A VGND VGND VPWR VPWR _16352_/X sky130_fd_sc_hd__buf_2
X_13564_ _13564_/A _13563_/X VGND VGND VPWR VPWR _13564_/X sky130_fd_sc_hd__or2_4
XFILLER_125_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20807__A _20832_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15303_ _15314_/A _15301_/X HADDR[23] _15301_/X VGND VGND VPWR VPWR _15303_/X sky130_fd_sc_hd__a2bb2o_4
X_12515_ _12328_/Y _12515_/B VGND VGND VPWR VPWR _12515_/X sky130_fd_sc_hd__or2_4
X_19071_ _19071_/A VGND VGND VPWR VPWR _19071_/X sky130_fd_sc_hd__buf_2
XFILLER_8_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13495_ _24967_/Q _13488_/X _13494_/Y VGND VGND VPWR VPWR _13495_/X sky130_fd_sc_hd__o21a_4
X_16283_ _14910_/Y _16278_/X _15982_/X _16282_/X VGND VGND VPWR VPWR _16283_/X sky130_fd_sc_hd__a2bb2o_4
X_18022_ _18022_/A VGND VGND VPWR VPWR _18022_/X sky130_fd_sc_hd__buf_2
X_12446_ _12415_/B _12415_/D _12423_/A VGND VGND VPWR VPWR _12458_/A sky130_fd_sc_hd__or3_4
X_15234_ _13770_/A _13780_/B _13782_/B VGND VGND VPWR VPWR _15234_/X sky130_fd_sc_hd__or3_4
XFILLER_51_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12377_ _25092_/Q VGND VGND VPWR VPWR _12415_/B sky130_fd_sc_hd__inv_2
X_15165_ _15165_/A _15165_/B _15164_/X VGND VGND VPWR VPWR _15165_/X sky130_fd_sc_hd__and3_4
XFILLER_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14116_ _14108_/Y _14115_/X VGND VGND VPWR VPWR _14116_/X sky130_fd_sc_hd__or2_4
X_15096_ _15096_/A _15144_/A VGND VGND VPWR VPWR _15097_/C sky130_fd_sc_hd__or2_4
X_19973_ _21953_/B _19970_/X _19445_/A _19970_/X VGND VGND VPWR VPWR _23141_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21638__A _21638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18924_ _23517_/Q VGND VGND VPWR VPWR _18924_/Y sky130_fd_sc_hd__inv_2
X_14047_ _14047_/A _17197_/B VGND VGND VPWR VPWR _14048_/A sky130_fd_sc_hd__nor2_4
XFILLER_136_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22206__A1_N _11985_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21421__B1 _21292_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18855_ _18851_/Y _18854_/X _18764_/X _18854_/X VGND VGND VPWR VPWR _18855_/X sky130_fd_sc_hd__a2bb2o_4
X_17806_ _17806_/A VGND VGND VPWR VPWR _17955_/A sky130_fd_sc_hd__buf_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18786_ _18782_/Y _18785_/X _18764_/X _18785_/X VGND VGND VPWR VPWR _23566_/D sky130_fd_sc_hd__a2bb2o_4
X_15998_ _15997_/Y _15993_/X _15801_/X _15993_/X VGND VGND VPWR VPWR _24362_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15651__A1 _15421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22469__A _24482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24246__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22516__A3 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17737_ _17783_/A _17737_/B _17736_/X VGND VGND VPWR VPWR _17737_/X sky130_fd_sc_hd__and3_4
X_14949_ _15177_/A _24272_/Q _24671_/Q _14900_/Y VGND VGND VPWR VPWR _14949_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA_clkbuf_5_20_0_HCLK_A clkbuf_4_10_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12995__A _12925_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13662__B1 _11607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21724__B2 _16041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17668_ _13406_/A _17666_/Y _17655_/X _17667_/X VGND VGND VPWR VPWR _17668_/X sky130_fd_sc_hd__o22a_4
XFILLER_63_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19407_ _19406_/Y _19402_/X _19360_/X _19402_/X VGND VGND VPWR VPWR _23346_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16600__B1 _24137_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16619_ _15657_/X _16597_/X _16558_/X _24125_/Q _16590_/X VGND VGND VPWR VPWR _16619_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_50_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17599_ _16700_/X _17605_/B VGND VGND VPWR VPWR _17603_/B sky130_fd_sc_hd__or2_4
XFILLER_56_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22916__B _23008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19338_ _23370_/Q VGND VGND VPWR VPWR _19338_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11976__B1 _11631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23881__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_245_0_HCLK clkbuf_8_245_0_HCLK/A VGND VGND VPWR VPWR _24662_/CLK sky130_fd_sc_hd__clkbuf_1
X_19269_ _19268_/Y _19266_/X _19221_/X _19266_/X VGND VGND VPWR VPWR _19269_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21300_ _21300_/A _21300_/B VGND VGND VPWR VPWR _21300_/Y sky130_fd_sc_hd__nor2_4
X_22280_ _22279_/X VGND VGND VPWR VPWR _22280_/X sky130_fd_sc_hd__buf_2
XANTENNA__12551__A2_N _24527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25034__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21231_ _14486_/X VGND VGND VPWR VPWR _21231_/X sky130_fd_sc_hd__buf_2
XANTENNA__12880__D _12854_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16667__B1 _16373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21162_ _21155_/X _21160_/X _21930_/A VGND VGND VPWR VPWR _21162_/X sky130_fd_sc_hd__o21a_4
X_20113_ _20112_/Y _20110_/X _19617_/A _20110_/X VGND VGND VPWR VPWR _20113_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14142__B2 _13492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21093_ _14936_/Y _21093_/B VGND VGND VPWR VPWR _21093_/X sky130_fd_sc_hd__and2_4
XFILLER_59_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16419__B1 _16254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21412__B1 _25193_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20044_ _20043_/Y _20041_/X _19721_/X _20041_/X VGND VGND VPWR VPWR _23114_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24921_ _24923_/CLK _13694_/X HRESETn VGND VGND VPWR VPWR _20402_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_28_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21963__A1 _21214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24852_ _24968_/CLK _24852_/D HRESETn VGND VGND VPWR VPWR _24852_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22379__A _21245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21283__A _21867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23803_ _23353_/CLK _23803_/D HRESETn VGND VGND VPWR VPWR _11706_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_22_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21995_ _22992_/B VGND VGND VPWR VPWR _21995_/X sky130_fd_sc_hd__buf_2
XANTENNA__13653__B1 _11590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24783_ _24783_/CLK _24783_/D HRESETn VGND VGND VPWR VPWR _23617_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20946_ _17646_/A VGND VGND VPWR VPWR _20946_/X sky130_fd_sc_hd__buf_2
XPHY_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23734_ _23734_/CLK _20589_/Y HRESETn VGND VGND VPWR VPWR _13533_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23969__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ _18632_/Y _17222_/B _21079_/B _20876_/Y VGND VGND VPWR VPWR _20878_/B sky130_fd_sc_hd__o22a_4
Xclkbuf_6_55_0_HCLK clkbuf_6_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_55_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23665_ _23661_/CLK _23665_/D HRESETn VGND VGND VPWR VPWR _23665_/Q sky130_fd_sc_hd__dfstp_4
XPHY_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22616_ _22616_/A VGND VGND VPWR VPWR _22616_/X sky130_fd_sc_hd__buf_2
XPHY_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23596_ _23596_/CLK _18698_/X VGND VGND VPWR VPWR _23596_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_70_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22140__A1 _11904_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11967__B1 _11612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19732__A2_N _19727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22547_ _22547_/A VGND VGND VPWR VPWR _22547_/X sky130_fd_sc_hd__buf_2
XANTENNA__20151__B1 _19963_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12300_ _12300_/A _12300_/B _12300_/C VGND VGND VPWR VPWR _12300_/X sky130_fd_sc_hd__and3_4
X_13280_ _13092_/A _19389_/A VGND VGND VPWR VPWR _13280_/X sky130_fd_sc_hd__or2_4
XFILLER_6_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22478_ _22226_/X _22477_/Y _16594_/Y _22228_/X VGND VGND VPWR VPWR _22478_/X sky130_fd_sc_hd__o22a_4
X_12231_ _12230_/X VGND VGND VPWR VPWR _12232_/B sky130_fd_sc_hd__inv_2
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21429_ _21066_/B VGND VGND VPWR VPWR _21434_/A sky130_fd_sc_hd__buf_2
X_24217_ _23840_/CLK _16407_/X HRESETn VGND VGND VPWR VPWR _24217_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22005__A2_N _22230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25197_ _23957_/CLK _11613_/X HRESETn VGND VGND VPWR VPWR _25197_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12392__B1 _12391_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12162_ _12120_/X _12162_/B VGND VGND VPWR VPWR _12502_/A sky130_fd_sc_hd__or2_4
X_24148_ _24113_/CLK _16582_/X HRESETn VGND VGND VPWR VPWR _24148_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24757__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15456__A _15455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12093_ _12084_/X _12093_/B _12090_/X _12092_/X VGND VGND VPWR VPWR _12093_/X sky130_fd_sc_hd__or4_4
X_16970_ _24310_/Q _16968_/Y _24316_/Q _17070_/A VGND VGND VPWR VPWR _16972_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15330__B1 _11525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24079_ _24079_/CLK _16892_/Y HRESETn VGND VGND VPWR VPWR _24079_/Q sky130_fd_sc_hd__dfrtp_4
X_15921_ _15921_/A VGND VGND VPWR VPWR _15921_/X sky130_fd_sc_hd__buf_2
XFILLER_1_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18640_ _23614_/Q VGND VGND VPWR VPWR _22056_/B sky130_fd_sc_hd__inv_2
XFILLER_7_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15852_ _15851_/Y _15847_/X _15765_/X _15847_/X VGND VGND VPWR VPWR _24417_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14803_ _24710_/Q VGND VGND VPWR VPWR _14882_/A sky130_fd_sc_hd__inv_2
X_18571_ _18571_/A _18568_/X _18569_/X _18571_/D VGND VGND VPWR VPWR _18571_/X sky130_fd_sc_hd__or4_4
X_15783_ _15781_/X _15763_/X _15499_/X _22420_/A _15779_/X VGND VGND VPWR VPWR _24443_/D
+ sky130_fd_sc_hd__a32o_4
X_12995_ _12925_/X _12974_/B _12994_/X VGND VGND VPWR VPWR _25010_/D sky130_fd_sc_hd__and3_4
X_17522_ _17521_/X VGND VGND VPWR VPWR _17522_/Y sky130_fd_sc_hd__inv_2
X_14734_ _14734_/A _14727_/X _14734_/C _14734_/D VGND VGND VPWR VPWR _14734_/X sky130_fd_sc_hd__or4_4
X_11946_ _11507_/X VGND VGND VPWR VPWR _15414_/A sky130_fd_sc_hd__buf_2
X_17453_ _17453_/A VGND VGND VPWR VPWR _17453_/X sky130_fd_sc_hd__buf_2
XFILLER_33_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15397__B1 _15279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21921__A _20975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14665_ _14665_/A VGND VGND VPWR VPWR _14665_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11877_ _11873_/X VGND VGND VPWR VPWR _11877_/Y sky130_fd_sc_hd__inv_2
X_16404_ _24218_/Q VGND VGND VPWR VPWR _16404_/Y sky130_fd_sc_hd__inv_2
X_13616_ _21293_/B VGND VGND VPWR VPWR _22439_/B sky130_fd_sc_hd__buf_2
XANTENNA__23639__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17384_ _17251_/Y _17382_/X _17383_/Y VGND VGND VPWR VPWR _17384_/X sky130_fd_sc_hd__o21a_4
X_14596_ _14596_/A VGND VGND VPWR VPWR _19189_/B sky130_fd_sc_hd__buf_2
XFILLER_32_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11958__B1 _11643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19123_ _14581_/Y _19123_/B _14587_/X _19123_/D VGND VGND VPWR VPWR _19123_/X sky130_fd_sc_hd__or4_4
XFILLER_9_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16335_ _16332_/Y _16333_/X _16334_/X _16333_/X VGND VGND VPWR VPWR _24243_/D sky130_fd_sc_hd__a2bb2o_4
X_13547_ _24964_/Q _13545_/X _13546_/Y VGND VGND VPWR VPWR _13547_/X sky130_fd_sc_hd__o21a_4
XANTENNA__20142__B1 _13668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22682__A2 _22011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19054_ _19053_/Y _19049_/X _18964_/X _19034_/Y VGND VGND VPWR VPWR _19054_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16266_ HWDATA[17] VGND VGND VPWR VPWR _16266_/X sky130_fd_sc_hd__buf_2
X_13478_ _13478_/A VGND VGND VPWR VPWR _13478_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_12_0_HCLK clkbuf_7_6_0_HCLK/X VGND VGND VPWR VPWR _23343_/CLK sky130_fd_sc_hd__clkbuf_1
X_18005_ _18005_/A VGND VGND VPWR VPWR _18005_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17268__D _17267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15217_ _15197_/X VGND VGND VPWR VPWR _15218_/B sky130_fd_sc_hd__inv_2
X_12429_ _12429_/A VGND VGND VPWR VPWR _12429_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_75_0_HCLK clkbuf_8_75_0_HCLK/A VGND VGND VPWR VPWR _25159_/CLK sky130_fd_sc_hd__clkbuf_1
X_16197_ _16195_/Y _16191_/X _15978_/X _16196_/X VGND VGND VPWR VPWR _24298_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15148_ _15138_/A _15146_/X _15147_/X VGND VGND VPWR VPWR _15148_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__21368__A _21235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24498__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15366__A _15358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24975__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15079_ _15057_/X _15079_/B _15078_/Y VGND VGND VPWR VPWR _24688_/D sky130_fd_sc_hd__and3_4
X_19956_ _19955_/Y _19953_/X _19381_/X _19953_/X VGND VGND VPWR VPWR _19956_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24427__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18907_ _18905_/Y _18900_/X _18883_/X _18906_/X VGND VGND VPWR VPWR _18907_/X sky130_fd_sc_hd__a2bb2o_4
X_19887_ _19887_/A VGND VGND VPWR VPWR _21960_/B sky130_fd_sc_hd__inv_2
XFILLER_67_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18838_ _18832_/Y VGND VGND VPWR VPWR _18838_/X sky130_fd_sc_hd__buf_2
XFILLER_68_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24080__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18769_ _18776_/A VGND VGND VPWR VPWR _18769_/X sky130_fd_sc_hd__buf_2
XFILLER_83_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20800_ _20800_/A VGND VGND VPWR VPWR _20800_/X sky130_fd_sc_hd__buf_2
X_21780_ _21777_/A _21780_/B VGND VGND VPWR VPWR _21780_/X sky130_fd_sc_hd__or2_4
XFILLER_51_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20731_ _23662_/Q VGND VGND VPWR VPWR _20733_/B sky130_fd_sc_hd__inv_2
XFILLER_63_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15388__B1 _15386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22713__A1_N _12410_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20920__A2 _20916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23450_ _23482_/CLK _19112_/X VGND VGND VPWR VPWR _17845_/B sky130_fd_sc_hd__dfxtp_4
X_20662_ _20647_/X _20661_/Y _16495_/A _20651_/X VGND VGND VPWR VPWR _20662_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25215__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22401_ _22401_/A _22265_/B VGND VGND VPWR VPWR _22401_/X sky130_fd_sc_hd__and2_4
X_23381_ _23374_/CLK _19309_/X VGND VGND VPWR VPWR _23381_/Q sky130_fd_sc_hd__dfxtp_4
X_20593_ _20592_/X VGND VGND VPWR VPWR _23735_/D sky130_fd_sc_hd__inv_2
XANTENNA__12610__B2 _24517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22332_ _22306_/X _22310_/X _22317_/Y _22331_/X VGND VGND VPWR VPWR HRDATA[11] sky130_fd_sc_hd__a211o_4
XANTENNA__20684__A1 _24996_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25120_ _25123_/CLK _25120_/D HRESETn VGND VGND VPWR VPWR _12116_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_104_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25051_ _24521_/CLK _12725_/Y HRESETn VGND VGND VPWR VPWR _12600_/A sky130_fd_sc_hd__dfrtp_4
X_22263_ _22223_/A VGND VGND VPWR VPWR _22263_/X sky130_fd_sc_hd__buf_2
XFILLER_136_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17756__A _14577_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19826__B1 _19825_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24002_ _25217_/CLK _17362_/X HRESETn VGND VGND VPWR VPWR _24002_/Q sky130_fd_sc_hd__dfrtp_4
X_21214_ _21214_/A _18659_/Y VGND VGND VPWR VPWR _21214_/X sky130_fd_sc_hd__or2_4
XFILLER_65_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22976__A3 _22839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22194_ _22193_/X VGND VGND VPWR VPWR _22194_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24850__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21145_ _21335_/A _21145_/B VGND VGND VPWR VPWR _21145_/X sky130_fd_sc_hd__or2_4
XANTENNA__15312__B1 HADDR[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22189__A1 _22444_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24168__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22189__B2 _22188_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21076_ _14282_/Y _20863_/A _23618_/Q _15639_/X VGND VGND VPWR VPWR _21076_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17065__B1 _17057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20027_ _20014_/Y VGND VGND VPWR VPWR _20027_/X sky130_fd_sc_hd__buf_2
X_24904_ _24904_/CLK _13909_/X HRESETn VGND VGND VPWR VPWR _24904_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23643__D scl_i_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24835_ _24851_/CLK _14162_/X HRESETn VGND VGND VPWR VPWR _24835_/Q sky130_fd_sc_hd__dfrtp_4
X_11800_ _11809_/A _17448_/B VGND VGND VPWR VPWR _11802_/A sky130_fd_sc_hd__or2_4
XFILLER_92_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12780_ _25011_/Q _12778_/Y _12779_/Y _22891_/A VGND VGND VPWR VPWR _12780_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24766_ _24851_/CLK _14396_/X HRESETn VGND VGND VPWR VPWR _13449_/A sky130_fd_sc_hd__dfrtp_4
X_21978_ _22527_/B VGND VGND VPWR VPWR _21978_/X sky130_fd_sc_hd__buf_2
XFILLER_15_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11731_ _23890_/Q VGND VGND VPWR VPWR _11732_/B sky130_fd_sc_hd__buf_2
XANTENNA__15379__B1 _13658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23717_ _23753_/CLK _23717_/D HRESETn VGND VGND VPWR VPWR _23717_/Q sky130_fd_sc_hd__dfrtp_4
X_20929_ _15405_/Y _22488_/B VGND VGND VPWR VPWR _20929_/X sky130_fd_sc_hd__and2_4
XPHY_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24697_ _24706_/CLK _15046_/X HRESETn VGND VGND VPWR VPWR _15044_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_14_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14450_ _21008_/A VGND VGND VPWR VPWR _21657_/A sky130_fd_sc_hd__buf_2
XFILLER_41_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23732__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _13591_/A _23917_/Q _13591_/A _23917_/Q VGND VGND VPWR VPWR _11669_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23648_ _23648_/CLK _20704_/X HRESETn VGND VGND VPWR VPWR _13998_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_30_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14051__B1 _13665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _20883_/A _13397_/Y _13330_/X _13397_/Y VGND VGND VPWR VPWR _24973_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11593_ HWDATA[12] VGND VGND VPWR VPWR _16096_/A sky130_fd_sc_hd__buf_2
X_14381_ _13435_/Y _14380_/X VGND VGND VPWR VPWR _14382_/B sky130_fd_sc_hd__or2_4
XANTENNA__20124__B1 _15520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22664__A2 _22662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12601__B2 _24516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23579_ _23563_/CLK _18748_/X VGND VGND VPWR VPWR _23579_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16120_ _16119_/Y _16117_/X _15282_/X _16117_/X VGND VGND VPWR VPWR _16120_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13332_ _13332_/A VGND VGND VPWR VPWR _13332_/Y sky130_fd_sc_hd__inv_2
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24938__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16051_ _16083_/A VGND VGND VPWR VPWR _16071_/A sky130_fd_sc_hd__buf_2
XANTENNA__14354__A1 scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13263_ _13159_/X _13261_/X _13263_/C VGND VGND VPWR VPWR _13264_/C sky130_fd_sc_hd__and3_4
X_15002_ _15001_/X VGND VGND VPWR VPWR _24708_/D sky130_fd_sc_hd__inv_2
X_12214_ _12538_/B _12214_/B _12213_/X VGND VGND VPWR VPWR _12215_/A sky130_fd_sc_hd__or3_4
XANTENNA__21188__A _21188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13194_ _11732_/B _13194_/B VGND VGND VPWR VPWR _13194_/X sky130_fd_sc_hd__or2_4
XANTENNA__22967__A3 _22251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24591__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12145_ _12180_/B _24549_/Q _25130_/Q _12144_/Y VGND VGND VPWR VPWR _12151_/B sky130_fd_sc_hd__a2bb2o_4
X_19810_ _19801_/A _18067_/A _13398_/A _13269_/B _19802_/A VGND VGND VPWR VPWR _23200_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_124_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15186__A _15158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15303__B1 HADDR[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24520__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12076_ _25129_/Q VGND VGND VPWR VPWR _12185_/A sky130_fd_sc_hd__inv_2
X_16953_ _16953_/A _16952_/Y _16951_/C VGND VGND VPWR VPWR _16953_/X sky130_fd_sc_hd__and3_4
X_19741_ _21925_/B _19738_/X _19714_/X _19738_/X VGND VGND VPWR VPWR _19741_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20820__A _20819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15904_ _24397_/Q VGND VGND VPWR VPWR _15904_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19672_ _23252_/Q VGND VGND VPWR VPWR _19672_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16884_ _16920_/A _16840_/B VGND VGND VPWR VPWR _16885_/B sky130_fd_sc_hd__or2_4
XFILLER_37_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18623_ _18622_/X VGND VGND VPWR VPWR _18624_/A sky130_fd_sc_hd__buf_2
XFILLER_77_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11652__A2_N _23914_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15835_ _15832_/Y _15827_/X _15753_/X _15834_/X VGND VGND VPWR VPWR _15835_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13434__A _24932_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18554_ _18422_/Y _18552_/X _18553_/Y VGND VGND VPWR VPWR _18554_/X sky130_fd_sc_hd__o21a_4
X_15766_ _12853_/Y _15757_/X _15765_/X _15757_/X VGND VGND VPWR VPWR _24451_/D sky130_fd_sc_hd__a2bb2o_4
X_12978_ _12992_/A _12976_/X _12977_/X VGND VGND VPWR VPWR _25016_/D sky130_fd_sc_hd__and3_4
XFILLER_46_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17505_ _17478_/Y _17505_/B _17505_/C _17505_/D VGND VGND VPWR VPWR _17505_/X sky130_fd_sc_hd__or4_4
X_14717_ _14716_/Y VGND VGND VPWR VPWR _15085_/A sky130_fd_sc_hd__buf_2
XANTENNA__21651__A _15824_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11929_ _11928_/Y _11924_/X _11930_/A _11924_/X VGND VGND VPWR VPWR _25160_/D sky130_fd_sc_hd__a2bb2o_4
X_18485_ _18518_/A _18515_/A _18485_/C _18485_/D VGND VGND VPWR VPWR _18507_/B sky130_fd_sc_hd__or4_4
X_15697_ _12346_/Y _15695_/X _15511_/X _15695_/X VGND VGND VPWR VPWR _15697_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22466__B _22246_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17436_ _17320_/A _17435_/X VGND VGND VPWR VPWR _17438_/A sky130_fd_sc_hd__nand2_4
X_14648_ _14621_/X _14646_/X _24629_/Q _14647_/X VGND VGND VPWR VPWR _14648_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__14042__B1 _13645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18308__B1 _18228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17367_ _17327_/D _17366_/X _17288_/Y VGND VGND VPWR VPWR _17368_/C sky130_fd_sc_hd__o21a_4
X_14579_ _17694_/A VGND VGND VPWR VPWR _17698_/A sky130_fd_sc_hd__buf_2
XANTENNA__15790__B1 _15511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19106_ _19114_/A VGND VGND VPWR VPWR _19106_/X sky130_fd_sc_hd__buf_2
XFILLER_105_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16318_ _24249_/Q VGND VGND VPWR VPWR _16318_/Y sky130_fd_sc_hd__inv_2
X_17298_ _17586_/A VGND VGND VPWR VPWR _17510_/B sky130_fd_sc_hd__buf_2
XANTENNA__22482__A _22263_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19037_ _13097_/B VGND VGND VPWR VPWR _19037_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24679__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16249_ _16228_/X _16234_/X _15477_/X _24281_/Q _16237_/X VGND VGND VPWR VPWR _16249_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16480__A _16530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24608__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13609__A _13460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16637__A3 HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24261__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19939_ _19926_/Y VGND VGND VPWR VPWR _19939_/X sky130_fd_sc_hd__buf_2
XFILLER_25_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15824__A _15824_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22950_ _22547_/X _22948_/X _22551_/X _22949_/X VGND VGND VPWR VPWR _22951_/B sky130_fd_sc_hd__o22a_4
XFILLER_96_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21901_ _24920_/Q _21720_/B VGND VGND VPWR VPWR _21905_/A sky130_fd_sc_hd__and2_4
X_22881_ _16056_/A _22549_/A _22864_/X VGND VGND VPWR VPWR _22881_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13344__A _13338_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_120_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_241_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24620_ _24620_/CLK _15306_/X HRESETn VGND VGND VPWR VPWR _24620_/Q sky130_fd_sc_hd__dfrtp_4
X_21832_ _20979_/A _21832_/B VGND VGND VPWR VPWR _21832_/X sky130_fd_sc_hd__or2_4
XFILLER_58_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14281__B1 _14213_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21736__A2_N _21083_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22657__A _21069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21561__A _22279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21763_ _21762_/X _21763_/B VGND VGND VPWR VPWR _21763_/X sky130_fd_sc_hd__or2_4
XFILLER_19_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24551_ _24566_/CLK _24551_/D HRESETn VGND VGND VPWR VPWR _12075_/A sky130_fd_sc_hd__dfrtp_4
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20714_ _23622_/Q _23623_/Q _20713_/Y VGND VGND VPWR VPWR _20714_/X sky130_fd_sc_hd__o21a_4
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23502_ _23537_/CLK _18971_/X VGND VGND VPWR VPWR _13041_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_51_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21694_ _22870_/B VGND VGND VPWR VPWR _21694_/X sky130_fd_sc_hd__buf_2
XANTENNA__14033__B1 _13668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24482_ _24478_/CLK _15687_/X HRESETn VGND VGND VPWR VPWR _24482_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20645_ _13524_/B _20639_/A _20644_/X VGND VGND VPWR VPWR _20645_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23433_ _23425_/CLK _23433_/D VGND VGND VPWR VPWR _17884_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_32_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23364_ _23350_/CLK _19356_/X VGND VGND VPWR VPWR _13137_/B sky130_fd_sc_hd__dfxtp_4
X_20576_ _20575_/Y _20570_/Y _13532_/B VGND VGND VPWR VPWR _20576_/X sky130_fd_sc_hd__o21a_4
XANTENNA__13510__C _13509_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20121__A3 _13668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25103_ _25115_/CLK _12300_/X HRESETn VGND VGND VPWR VPWR _12299_/A sky130_fd_sc_hd__dfrtp_4
X_22315_ _22264_/X _22314_/X _16358_/Y _16305_/X VGND VGND VPWR VPWR _22315_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23295_ _23383_/CLK _23295_/D VGND VGND VPWR VPWR _23295_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16390__A _11527_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12347__B1 _12345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24349__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22246_ _16193_/A _22246_/B VGND VGND VPWR VPWR _22246_/X sky130_fd_sc_hd__or2_4
X_25034_ _25034_/CLK _25034_/D HRESETn VGND VGND VPWR VPWR _12812_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_79_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22177_ _11606_/Y _22857_/B _15981_/A _16134_/X VGND VGND VPWR VPWR _22177_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21128_ _21071_/X _21091_/X _21128_/C _21127_/X VGND VGND VPWR VPWR _21128_/X sky130_fd_sc_hd__or4_4
XFILLER_121_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13950_ _13950_/A _13937_/A VGND VGND VPWR VPWR _13950_/X sky130_fd_sc_hd__and2_4
X_21059_ _22933_/B VGND VGND VPWR VPWR _21059_/X sky130_fd_sc_hd__buf_2
XFILLER_47_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18786__B1 _18764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22582__A1 _16078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12901_ _12812_/A _12900_/Y VGND VGND VPWR VPWR _12901_/X sky130_fd_sc_hd__or2_4
XANTENNA__23984__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13881_ _13881_/A VGND VGND VPWR VPWR _13898_/A sky130_fd_sc_hd__inv_2
XANTENNA__16683__A2_N _22307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15620_ _15619_/X _15617_/X _15507_/X _24513_/Q _15585_/A VGND VGND VPWR VPWR _24513_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_59_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12832_ _22419_/A VGND VGND VPWR VPWR _12880_/B sky130_fd_sc_hd__inv_2
XFILLER_34_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23913__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24818_ _24788_/CLK _24818_/D HRESETn VGND VGND VPWR VPWR _21073_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25137__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22567__A _22681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15551_ _15549_/Y _15546_/X _15550_/X _15546_/X VGND VGND VPWR VPWR _24538_/D sky130_fd_sc_hd__a2bb2o_4
X_12763_ _12584_/Y _12762_/X VGND VGND VPWR VPWR _12765_/B sky130_fd_sc_hd__or2_4
XPHY_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24749_ _24748_/CLK _14516_/X HRESETn VGND VGND VPWR VPWR _24749_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16565__A _22228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _21751_/A VGND VGND VPWR VPWR _14502_/Y sky130_fd_sc_hd__inv_2
XPHY_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11697_/Y _11711_/X VGND VGND VPWR VPWR _11714_/X sky130_fd_sc_hd__and2_4
X_18270_ _18207_/B _18265_/B _18237_/X _18266_/Y VGND VGND VPWR VPWR _18270_/X sky130_fd_sc_hd__a211o_4
XFILLER_37_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _11532_/X VGND VGND VPWR VPWR _15482_/X sky130_fd_sc_hd__buf_2
XPHY_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12637_/X _12694_/B _12693_/X VGND VGND VPWR VPWR _25060_/D sky130_fd_sc_hd__and3_4
XPHY_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_25_0_HCLK clkbuf_4_12_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _17220_/X VGND VGND VPWR VPWR _17222_/B sky130_fd_sc_hd__buf_2
XPHY_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14433_/A _14432_/X VGND VGND VPWR VPWR _14433_/X sky130_fd_sc_hd__and2_4
XFILLER_52_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _23802_/Q VGND VGND VPWR VPWR _11645_/X sky130_fd_sc_hd__buf_2
XANTENNA__19876__A _19876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17152_ _17034_/C _17134_/X VGND VGND VPWR VPWR _17152_/Y sky130_fd_sc_hd__nand2_4
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14364_ _24769_/Q _13893_/X _13887_/X VGND VGND VPWR VPWR _24769_/D sky130_fd_sc_hd__a21bo_4
X_11576_ HWDATA[16] VGND VGND VPWR VPWR _11576_/X sky130_fd_sc_hd__buf_2
XFILLER_11_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20815__A _20814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16103_ _22267_/A _16099_/X _15788_/X _16099_/X VGND VGND VPWR VPWR _16103_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24772__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13315_ _13219_/A _23335_/Q VGND VGND VPWR VPWR _13315_/X sky130_fd_sc_hd__or2_4
X_17083_ _17074_/A VGND VGND VPWR VPWR _17083_/X sky130_fd_sc_hd__buf_2
XFILLER_122_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15524__B1 _15286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14295_ _24788_/Q VGND VGND VPWR VPWR _14295_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24701__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16034_ _19144_/B _16033_/B _16032_/Y _16033_/Y VGND VGND VPWR VPWR _16034_/X sky130_fd_sc_hd__a211o_4
X_13246_ _13278_/A _13244_/X _13245_/X VGND VGND VPWR VPWR _13246_/X sky130_fd_sc_hd__and3_4
XANTENNA__19805__A3 _13668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24019__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16619__A3 _16558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13177_ _13244_/A _23475_/Q VGND VGND VPWR VPWR _13177_/X sky130_fd_sc_hd__or2_4
XFILLER_111_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11561__A1 _11533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_149_0_HCLK clkbuf_7_74_0_HCLK/X VGND VGND VPWR VPWR _24385_/CLK sky130_fd_sc_hd__clkbuf_1
X_12128_ _12127_/Y _24557_/Q _12127_/Y _24557_/Q VGND VGND VPWR VPWR _12131_/C sky130_fd_sc_hd__a2bb2o_4
X_17985_ _11691_/Y _17977_/X _15501_/X _17977_/X VGND VGND VPWR VPWR _23923_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20550__A _20550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12059_ _25135_/Q VGND VGND VPWR VPWR SSn_S3 sky130_fd_sc_hd__inv_2
X_16936_ _16936_/A _16936_/B _16935_/Y VGND VGND VPWR VPWR _16936_/X sky130_fd_sc_hd__and3_4
X_19724_ _19724_/A VGND VGND VPWR VPWR _19724_/X sky130_fd_sc_hd__buf_2
XFILLER_78_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16867_ _16867_/A _16867_/B _16866_/X VGND VGND VPWR VPWR _16867_/X sky130_fd_sc_hd__and3_4
X_19655_ _19654_/Y _19652_/X _19607_/X _19652_/X VGND VGND VPWR VPWR _23259_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13164__A _13073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15818_ _24426_/Q VGND VGND VPWR VPWR _15818_/Y sky130_fd_sc_hd__inv_2
X_18606_ _23642_/Q VGND VGND VPWR VPWR _18607_/A sky130_fd_sc_hd__inv_2
XANTENNA__23654__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19586_ _21514_/B _19581_/X _19455_/X _19581_/X VGND VGND VPWR VPWR _19586_/X sky130_fd_sc_hd__a2bb2o_4
X_16798_ _16798_/A VGND VGND VPWR VPWR _16853_/A sky130_fd_sc_hd__inv_2
XFILLER_53_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14263__B1 _14094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22325__A1 _22322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22477__A _22477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18537_ _18532_/A _18536_/X _18449_/X VGND VGND VPWR VPWR _18537_/Y sky130_fd_sc_hd__a21oi_4
X_15749_ _15748_/X _15740_/X _15468_/X _24459_/Q _15746_/X VGND VGND VPWR VPWR _24459_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_34_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22196__B _20757_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18468_ _18468_/A _18468_/B _18468_/C VGND VGND VPWR VPWR _18468_/X sky130_fd_sc_hd__or3_4
X_17419_ _17423_/A _17419_/B _17418_/Y VGND VGND VPWR VPWR _23988_/D sky130_fd_sc_hd__and3_4
X_18399_ _23835_/Q VGND VGND VPWR VPWR _18468_/A sky130_fd_sc_hd__inv_2
XANTENNA__12508__A _12508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22924__B _22857_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20430_ _20429_/Y _13500_/X _13503_/B VGND VGND VPWR VPWR _20430_/X sky130_fd_sc_hd__o21a_4
XFILLER_105_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18701__B1 _18700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20361_ _14052_/Y _20344_/X _20358_/X _20360_/X VGND VGND VPWR VPWR _20361_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15515__B1 _15513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15819__A _11529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22100_ _20961_/A _22100_/B VGND VGND VPWR VPWR _22100_/X sky130_fd_sc_hd__or2_4
XANTENNA__24442__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23080_ _23109_/CLK _23080_/D VGND VGND VPWR VPWR _23080_/Q sky130_fd_sc_hd__dfxtp_4
X_20292_ _20292_/A _20289_/A VGND VGND VPWR VPWR _20292_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_7_45_0_HCLK clkbuf_7_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_91_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15530__A3 _15432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22031_ _18110_/Y _20800_/A VGND VGND VPWR VPWR _22031_/X sky130_fd_sc_hd__and2_4
XANTENNA__13339__A _13338_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20811__A1 _24545_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15554__A _19452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22013__B1 _21867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23982_ _23990_/CLK _17433_/Y HRESETn VGND VGND VPWR VPWR _23982_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22933_ _16485_/Y _22933_/B VGND VGND VPWR VPWR _22933_/X sky130_fd_sc_hd__and2_4
XANTENNA__13074__A _13271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22864_ _22351_/A VGND VGND VPWR VPWR _22864_/X sky130_fd_sc_hd__buf_2
XANTENNA__15597__A3 _15596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14254__B1 _14236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24603_ _23744_/CLK _15356_/X HRESETn VGND VGND VPWR VPWR _24603_/Q sky130_fd_sc_hd__dfrtp_4
X_21815_ _20964_/A _20081_/Y VGND VGND VPWR VPWR _21815_/X sky130_fd_sc_hd__or2_4
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22795_ _15846_/Y _21042_/A _16157_/Y _21543_/A VGND VGND VPWR VPWR _22795_/X sky130_fd_sc_hd__o22a_4
XFILLER_24_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24534_ _25061_/CLK _15567_/X HRESETn VGND VGND VPWR VPWR _19859_/A sky130_fd_sc_hd__dfrtp_4
X_21746_ _21746_/A _15639_/X VGND VGND VPWR VPWR _21746_/X sky130_fd_sc_hd__and2_4
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15754__B1 _15753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24465_ _23442_/CLK _15732_/X HRESETn VGND VGND VPWR VPWR _24465_/Q sky130_fd_sc_hd__dfrtp_4
X_21677_ _21677_/A _21677_/B VGND VGND VPWR VPWR _21678_/C sky130_fd_sc_hd__or2_4
XANTENNA__12418__A _12391_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23416_ _23416_/CLK _23416_/D VGND VGND VPWR VPWR _19206_/A sky130_fd_sc_hd__dfxtp_4
X_20628_ _20635_/C _20653_/A _20627_/Y VGND VGND VPWR VPWR _20628_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24396_ _24399_/CLK _24396_/D HRESETn VGND VGND VPWR VPWR _24396_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15506__B1 _24557_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20559_ _13526_/A _13526_/B _13527_/B VGND VGND VPWR VPWR _20559_/Y sky130_fd_sc_hd__a21oi_4
X_23347_ _23336_/CLK _23347_/D VGND VGND VPWR VPWR _19404_/A sky130_fd_sc_hd__dfxtp_4
X_13100_ _13047_/A _13097_/X _13099_/X VGND VGND VPWR VPWR _13100_/X sky130_fd_sc_hd__and3_4
XFILLER_138_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24183__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14080_ _14077_/Y _14079_/X _13663_/X _14079_/X VGND VGND VPWR VPWR _14080_/X sky130_fd_sc_hd__a2bb2o_4
X_23278_ _23278_/CLK _23278_/D VGND VGND VPWR VPWR _23278_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15521__A3 _15520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24112__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13031_ _13047_/A _13028_/X _13030_/X VGND VGND VPWR VPWR _13031_/X sky130_fd_sc_hd__and3_4
XANTENNA__22252__B1 _24555_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25017_ _24451_/CLK _25017_/D HRESETn VGND VGND VPWR VPWR _22377_/A sky130_fd_sc_hd__dfrtp_4
X_22229_ _22226_/X _22227_/X _14821_/Y _22228_/X VGND VGND VPWR VPWR _22229_/X sky130_fd_sc_hd__o22a_4
XFILLER_65_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21466__A _21469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_2_0_HCLK clkbuf_6_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__15464__A _15463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17770_ _17916_/A _23452_/Q VGND VGND VPWR VPWR _17770_/X sky130_fd_sc_hd__or2_4
X_14982_ _14982_/A _15094_/A VGND VGND VPWR VPWR _14982_/X sky130_fd_sc_hd__and2_4
XFILLER_93_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16721_ _17489_/C VGND VGND VPWR VPWR _17614_/A sky130_fd_sc_hd__buf_2
X_13933_ _13933_/A _13931_/Y _13947_/A VGND VGND VPWR VPWR _13934_/C sky130_fd_sc_hd__and3_4
X_19440_ _19440_/A VGND VGND VPWR VPWR _19440_/Y sky130_fd_sc_hd__inv_2
X_16652_ _16624_/A VGND VGND VPWR VPWR _16652_/X sky130_fd_sc_hd__buf_2
X_13864_ _13852_/A _13828_/C _13880_/C VGND VGND VPWR VPWR _13864_/X sky130_fd_sc_hd__or3_4
XANTENNA__14245__B1 _14094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21185__A1_N _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22297__A _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15603_ _15588_/Y VGND VGND VPWR VPWR _15604_/A sky130_fd_sc_hd__buf_2
X_12815_ _22203_/A VGND VGND VPWR VPWR _12815_/Y sky130_fd_sc_hd__inv_2
X_19371_ _19799_/A _11761_/A _20134_/C VGND VGND VPWR VPWR _19372_/A sky130_fd_sc_hd__or3_4
X_16583_ _24147_/Q VGND VGND VPWR VPWR _16583_/Y sky130_fd_sc_hd__inv_2
X_13795_ _13795_/A VGND VGND VPWR VPWR _13796_/A sky130_fd_sc_hd__inv_2
X_18322_ _18322_/A _18322_/B VGND VGND VPWR VPWR _18323_/B sky130_fd_sc_hd__or2_4
X_15534_ _19442_/A VGND VGND VPWR VPWR _15534_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12746_ _12648_/Y _12742_/X VGND VGND VPWR VPWR _12746_/Y sky130_fd_sc_hd__nand2_4
XFILLER_72_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21530__A2 _21528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18253_ _18242_/B _18257_/B VGND VGND VPWR VPWR _18253_/Y sky130_fd_sc_hd__nand2_4
XFILLER_128_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24953__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15465_ _15464_/X VGND VGND VPWR VPWR _15466_/A sky130_fd_sc_hd__buf_2
XFILLER_124_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12677_ _12638_/Y _12653_/X _12612_/Y _12646_/X VGND VGND VPWR VPWR _12677_/X sky130_fd_sc_hd__or4_4
XANTENNA__12328__A _12328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ _24017_/Q VGND VGND VPWR VPWR _17204_/Y sky130_fd_sc_hd__inv_2
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ _14380_/B _14414_/X _14412_/X _14415_/X _14414_/A VGND VGND VPWR VPWR _24758_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_128_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11628_ _25193_/Q VGND VGND VPWR VPWR _11628_/Y sky130_fd_sc_hd__inv_2
X_18184_ _24346_/Q _18240_/C _16073_/Y _23865_/Q VGND VGND VPWR VPWR _18185_/D sky130_fd_sc_hd__a2bb2o_4
X_15396_ _15401_/A VGND VGND VPWR VPWR _15396_/X sky130_fd_sc_hd__buf_2
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15760__A3 _15596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17135_ _17034_/X _17134_/X VGND VGND VPWR VPWR _17135_/X sky130_fd_sc_hd__or2_4
X_14347_ _23649_/Q _14346_/X _14306_/A _14320_/Y VGND VGND VPWR VPWR _24772_/D sky130_fd_sc_hd__o22a_4
XFILLER_116_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22491__B1 _13509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11559_ _11541_/X VGND VGND VPWR VPWR _11559_/X sky130_fd_sc_hd__buf_2
XFILLER_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17066_ _17066_/A VGND VGND VPWR VPWR _17066_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14278_ _14277_/Y _14273_/X _14221_/X _14273_/X VGND VGND VPWR VPWR _24795_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23035__A2 _21703_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16017_ _16014_/A _16014_/B _16005_/X VGND VGND VPWR VPWR _16017_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_83_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13229_ _13261_/A _18981_/A VGND VGND VPWR VPWR _13231_/B sky130_fd_sc_hd__or2_4
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12063__A _12062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12998__A _12793_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15374__A _15358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23835__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17968_ _17968_/A _17968_/B _17967_/X VGND VGND VPWR VPWR _17968_/X sky130_fd_sc_hd__and3_4
XANTENNA__25059__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19707_ _23238_/Q VGND VGND VPWR VPWR _22091_/B sky130_fd_sc_hd__inv_2
X_16919_ _16919_/A VGND VGND VPWR VPWR _24071_/D sky130_fd_sc_hd__inv_2
X_17899_ _17899_/A _23529_/Q VGND VGND VPWR VPWR _17899_/X sky130_fd_sc_hd__or2_4
XANTENNA__18685__A _16216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19638_ _23264_/Q VGND VGND VPWR VPWR _21145_/B sky130_fd_sc_hd__inv_2
XFILLER_81_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19569_ _23288_/Q VGND VGND VPWR VPWR _21158_/B sky130_fd_sc_hd__inv_2
XANTENNA__22000__A _15456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21600_ _21585_/X _21600_/B _21600_/C _21599_/Y VGND VGND VPWR VPWR _21600_/X sky130_fd_sc_hd__and4_4
X_22580_ _24208_/Q _22580_/B VGND VGND VPWR VPWR _22580_/X sky130_fd_sc_hd__or2_4
XANTENNA__24694__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21531_ _23394_/Q _14016_/A _19223_/A _22042_/B VGND VGND VPWR VPWR _21531_/X sky130_fd_sc_hd__o22a_4
XFILLER_138_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24623__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21462_ _21169_/A _21462_/B VGND VGND VPWR VPWR _21464_/B sky130_fd_sc_hd__or2_4
X_24250_ _24225_/CLK _24250_/D HRESETn VGND VGND VPWR VPWR _24250_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20413_ _20413_/A VGND VGND VPWR VPWR _20414_/A sky130_fd_sc_hd__inv_2
XFILLER_135_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23201_ _24008_/CLK _23201_/D VGND VGND VPWR VPWR _23201_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15549__A _19452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21393_ _21393_/A _19830_/Y VGND VGND VPWR VPWR _21394_/C sky130_fd_sc_hd__or2_4
X_24181_ _24177_/CLK _16500_/X HRESETn VGND VGND VPWR VPWR _24181_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20344_ _20343_/Y VGND VGND VPWR VPWR _20344_/X sky130_fd_sc_hd__buf_2
X_23132_ _23133_/CLK _23132_/D VGND VGND VPWR VPWR _23132_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16161__B1 _15484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23063_ _20741_/X VGND VGND VPWR VPWR IRQ[11] sky130_fd_sc_hd__buf_2
X_20275_ _13996_/Y _20273_/X _14266_/X _20274_/X VGND VGND VPWR VPWR _20276_/A sky130_fd_sc_hd__a211o_4
XANTENNA__14711__B2 _22857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22014_ _22014_/A _22014_/B VGND VGND VPWR VPWR _22014_/X sky130_fd_sc_hd__and2_4
XFILLER_118_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_132_0_HCLK clkbuf_7_66_0_HCLK/X VGND VGND VPWR VPWR _23568_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_195_0_HCLK clkbuf_7_97_0_HCLK/X VGND VGND VPWR VPWR _24289_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13516__B _13515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23965_ _23969_/CLK _23965_/D HRESETn VGND VGND VPWR VPWR _17481_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22916_ _24495_/Q _23008_/B VGND VGND VPWR VPWR _22916_/X sky130_fd_sc_hd__or2_4
XFILLER_72_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21733__B _21716_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23896_ _23979_/CLK _18073_/X HRESETn VGND VGND VPWR VPWR _23896_/Q sky130_fd_sc_hd__dfrtp_4
X_22847_ _16475_/A VGND VGND VPWR VPWR _23020_/B sky130_fd_sc_hd__buf_2
XFILLER_71_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12600_ _12600_/A VGND VGND VPWR VPWR _12644_/D sky130_fd_sc_hd__inv_2
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13580_ _13580_/A VGND VGND VPWR VPWR _13580_/X sky130_fd_sc_hd__buf_2
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22778_ _22778_/A _11964_/A VGND VGND VPWR VPWR _22781_/B sky130_fd_sc_hd__or2_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12531_ _12534_/A _12537_/B VGND VGND VPWR VPWR _12535_/B sky130_fd_sc_hd__or2_4
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24517_ _24483_/CLK _24517_/D HRESETn VGND VGND VPWR VPWR _24517_/Q sky130_fd_sc_hd__dfrtp_4
X_21729_ _21729_/A _20832_/A VGND VGND VPWR VPWR _21729_/X sky130_fd_sc_hd__and2_4
XFILLER_38_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12148__A _24567_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22564__B _22564_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24364__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15250_ _15250_/A VGND VGND VPWR VPWR _15250_/X sky130_fd_sc_hd__buf_2
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12462_ _12444_/A _12458_/Y _12461_/X VGND VGND VPWR VPWR _12463_/A sky130_fd_sc_hd__or3_4
XFILLER_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24448_ _24445_/CLK _15774_/X HRESETn VGND VGND VPWR VPWR _22633_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_32_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15742__A3 _15735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14201_ _14201_/A VGND VGND VPWR VPWR _14201_/X sky130_fd_sc_hd__buf_2
XFILLER_138_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11987__A _11986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15181_ _15168_/X VGND VGND VPWR VPWR _15182_/B sky130_fd_sc_hd__inv_2
XFILLER_138_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15459__A _15459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12393_ _25098_/Q _12380_/Y _12379_/Y _21567_/A VGND VGND VPWR VPWR _12396_/C sky130_fd_sc_hd__a2bb2o_4
X_24379_ _24361_/CLK _15954_/X HRESETn VGND VGND VPWR VPWR _22639_/A sky130_fd_sc_hd__dfrtp_4
X_14132_ _14126_/X _14130_/X _13341_/A _14131_/X VGND VGND VPWR VPWR _24847_/D sky130_fd_sc_hd__o22a_4
XFILLER_67_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23017__A2 _22859_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14063_ _14062_/Y _14060_/X _13398_/X _14060_/X VGND VGND VPWR VPWR _14063_/X sky130_fd_sc_hd__a2bb2o_4
X_18940_ _17966_/B VGND VGND VPWR VPWR _18940_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13014_ _23890_/Q VGND VGND VPWR VPWR _13078_/A sky130_fd_sc_hd__inv_2
X_18871_ _18870_/Y _18866_/X _18828_/X _18854_/A VGND VGND VPWR VPWR _18871_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_91_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_91_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17822_ _17783_/A _17819_/X _17821_/X VGND VGND VPWR VPWR _17822_/X sky130_fd_sc_hd__and3_4
XFILLER_58_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25152__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22528__B2 _22121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14965_ _14964_/Y _24258_/Q _24651_/Q _14936_/Y VGND VGND VPWR VPWR _14965_/X sky130_fd_sc_hd__a2bb2o_4
X_17753_ _17918_/A VGND VGND VPWR VPWR _17961_/A sky130_fd_sc_hd__buf_2
XFILLER_48_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13916_ _13908_/A VGND VGND VPWR VPWR _13916_/X sky130_fd_sc_hd__buf_2
X_16704_ _16704_/A VGND VGND VPWR VPWR _17490_/B sky130_fd_sc_hd__inv_2
XFILLER_78_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17684_ _14573_/A _17684_/B VGND VGND VPWR VPWR _17684_/X sky130_fd_sc_hd__or2_4
XFILLER_63_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14896_ _15179_/A _24271_/Q _14895_/A _24271_/Q VGND VGND VPWR VPWR _14896_/X sky130_fd_sc_hd__a2bb2o_4
X_16635_ _16624_/X _16625_/X HWDATA[25] _24118_/Q _16622_/X VGND VGND VPWR VPWR _24118_/D
+ sky130_fd_sc_hd__a32o_4
X_19423_ _23340_/Q VGND VGND VPWR VPWR _19423_/Y sky130_fd_sc_hd__inv_2
X_13847_ _13845_/X _13846_/X VGND VGND VPWR VPWR _13847_/Y sky130_fd_sc_hd__nand2_4
XFILLER_50_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16566_ _16566_/A VGND VGND VPWR VPWR _16566_/X sky130_fd_sc_hd__buf_2
X_19354_ _13137_/B VGND VGND VPWR VPWR _19354_/Y sky130_fd_sc_hd__inv_2
X_13778_ _13778_/A VGND VGND VPWR VPWR _13779_/D sky130_fd_sc_hd__inv_2
XANTENNA__22755__A _22754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18904__B1 _18880_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15517_ _12075_/Y _15514_/X _15390_/X _15514_/X VGND VGND VPWR VPWR _24551_/D sky130_fd_sc_hd__a2bb2o_4
X_18305_ _18210_/B _18304_/X VGND VGND VPWR VPWR _18312_/B sky130_fd_sc_hd__or2_4
X_12729_ _12728_/X VGND VGND VPWR VPWR _12730_/B sky130_fd_sc_hd__inv_2
X_19285_ _22103_/B _19284_/X _11835_/X _19284_/X VGND VGND VPWR VPWR _23390_/D sky130_fd_sc_hd__a2bb2o_4
X_16497_ _24181_/Q VGND VGND VPWR VPWR _16497_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18236_ _18226_/A _18236_/B _18235_/X VGND VGND VPWR VPWR _18236_/X sky130_fd_sc_hd__and3_4
XFILLER_31_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15448_ _14433_/A _15447_/X _15445_/Y VGND VGND VPWR VPWR _24579_/D sky130_fd_sc_hd__o21a_4
XFILLER_50_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24034__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18167_ _18334_/A VGND VGND VPWR VPWR _18167_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22464__B1 _24517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15369__A HWDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15379_ _22278_/A _15374_/X _13658_/X _15374_/X VGND VGND VPWR VPWR _15379_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17118_ _24042_/Q _17117_/Y VGND VGND VPWR VPWR _17118_/X sky130_fd_sc_hd__or2_4
XFILLER_116_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18098_ _18089_/A _17226_/X _18097_/X VGND VGND VPWR VPWR _18099_/A sky130_fd_sc_hd__a21o_4
XANTENNA__22490__A _22407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17049_ _17048_/X VGND VGND VPWR VPWR _17051_/B sky130_fd_sc_hd__inv_2
X_20060_ _20060_/A VGND VGND VPWR VPWR _20060_/X sky130_fd_sc_hd__buf_2
XANTENNA__13617__A _22439_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_205_0_HCLK clkbuf_8_205_0_HCLK/A VGND VGND VPWR VPWR _24168_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15832__A _24424_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23750_ _24180_/CLK _23750_/D HRESETn VGND VGND VPWR VPWR _20656_/A sky130_fd_sc_hd__dfrtp_4
X_20962_ _20962_/A _20958_/X _20962_/C VGND VGND VPWR VPWR _20962_/X sky130_fd_sc_hd__and3_4
XANTENNA__24875__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22701_ _22195_/X _22700_/X _22629_/X _12088_/A _22198_/X VGND VGND VPWR VPWR _22702_/B
+ sky130_fd_sc_hd__a32o_4
X_23681_ _24769_/CLK scl_i_S5 HRESETn VGND VGND VPWR VPWR _23681_/Q sky130_fd_sc_hd__dfrtp_4
X_20893_ _11936_/Y _11954_/A _20892_/X VGND VGND VPWR VPWR _20893_/X sky130_fd_sc_hd__o21a_4
X_22632_ _21848_/B VGND VGND VPWR VPWR _22703_/B sky130_fd_sc_hd__buf_2
XFILLER_55_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17759__A _14571_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22563_ _20814_/X VGND VGND VPWR VPWR _22681_/A sky130_fd_sc_hd__buf_2
XANTENNA__16663__A _16643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24302_ _24031_/CLK _24302_/D HRESETn VGND VGND VPWR VPWR _16186_/A sky130_fd_sc_hd__dfrtp_4
X_21514_ _21383_/A _21514_/B VGND VGND VPWR VPWR _21515_/C sky130_fd_sc_hd__or2_4
XANTENNA__16382__B1 _16211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22494_ _22493_/X VGND VGND VPWR VPWR _22495_/D sky130_fd_sc_hd__inv_2
XFILLER_21_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21258__A1 _22146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24233_ _24201_/CLK _16360_/X HRESETn VGND VGND VPWR VPWR _16358_/A sky130_fd_sc_hd__dfrtp_4
X_21445_ _14257_/Y _11503_/A _14297_/A _15426_/X VGND VGND VPWR VPWR _21445_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19320__B1 _19227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21376_ _21376_/A _21374_/X _21375_/X VGND VGND VPWR VPWR _21376_/X sky130_fd_sc_hd__and3_4
X_24164_ _24167_/CLK _24164_/D HRESETn VGND VGND VPWR VPWR _16539_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_120_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20327_ _13955_/Y _20296_/A _20286_/X _20326_/Y VGND VGND VPWR VPWR _20328_/A sky130_fd_sc_hd__a211o_4
XANTENNA__17494__A _22376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23115_ _23939_/CLK _20042_/X VGND VGND VPWR VPWR _20040_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__23757__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21728__B _21425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24095_ _24101_/CLK _24095_/D HRESETn VGND VGND VPWR VPWR _14747_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22758__A1 _22195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_15_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_30_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_135_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22758__B2 _22198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20258_ _14099_/A _20243_/C _20257_/X VGND VGND VPWR VPWR _20265_/B sky130_fd_sc_hd__a21o_4
X_23046_ VGND VGND VPWR VPWR _23046_/HI IRQ[14] sky130_fd_sc_hd__conb_1
XANTENNA__20769__B1 _22884_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13650__A1_N _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20189_ _20189_/A _20189_/B VGND VGND VPWR VPWR _20194_/B sky130_fd_sc_hd__and2_4
XFILLER_88_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24997_ _23990_/CLK _24997_/D HRESETn VGND VGND VPWR VPWR _24997_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_92_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14750_ _14705_/X _14750_/B _14734_/X _14749_/X VGND VGND VPWR VPWR _14750_/X sky130_fd_sc_hd__or4_4
X_11962_ _11961_/X VGND VGND VPWR VPWR _22564_/B sky130_fd_sc_hd__buf_2
XFILLER_45_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_1_HCLK clkbuf_1_1_1_HCLK/A VGND VGND VPWR VPWR clkbuf_2_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_23948_ _23972_/CLK _17607_/X HRESETn VGND VGND VPWR VPWR _16685_/A sky130_fd_sc_hd__dfrtp_4
X_13701_ _13697_/X _13700_/X _24859_/Q _13693_/X VGND VGND VPWR VPWR _13701_/X sky130_fd_sc_hd__o22a_4
X_14681_ _14681_/A _14633_/A VGND VGND VPWR VPWR _14682_/A sky130_fd_sc_hd__or2_4
X_11893_ _24980_/Q _11881_/A _24980_/Q _11881_/A VGND VGND VPWR VPWR _11893_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16592__A1_N _14838_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23879_ _25141_/CLK _23879_/D HRESETn VGND VGND VPWR VPWR _18127_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16420_ _24211_/Q VGND VGND VPWR VPWR _16420_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24545__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13632_ _13632_/A VGND VGND VPWR VPWR _13632_/X sky130_fd_sc_hd__buf_2
XFILLER_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22575__A _22840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16351_ _24236_/Q VGND VGND VPWR VPWR _16351_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21497__A1 _21489_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13563_ _11673_/Y _13562_/X VGND VGND VPWR VPWR _13563_/X sky130_fd_sc_hd__or2_4
X_15302_ _11507_/A _15301_/X HWRITE _15301_/X VGND VGND VPWR VPWR _24623_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22294__B _22238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12514_ _12407_/B _12511_/D VGND VGND VPWR VPWR _12515_/B sky130_fd_sc_hd__or2_4
X_19070_ _17880_/B VGND VGND VPWR VPWR _19070_/Y sky130_fd_sc_hd__inv_2
X_16282_ _16262_/A VGND VGND VPWR VPWR _16282_/X sky130_fd_sc_hd__buf_2
X_13494_ _24967_/Q _13492_/X _13521_/A VGND VGND VPWR VPWR _13494_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_90_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18021_ _17625_/Y VGND VGND VPWR VPWR _18061_/B sky130_fd_sc_hd__buf_2
X_15233_ _15232_/X VGND VGND VPWR VPWR _24650_/D sky130_fd_sc_hd__inv_2
X_12445_ _12444_/X VGND VGND VPWR VPWR _25096_/D sky130_fd_sc_hd__inv_2
XANTENNA__22446__B1 _22435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14524__C _14521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15164_ _15104_/Y _15162_/A VGND VGND VPWR VPWR _15164_/X sky130_fd_sc_hd__or2_4
X_12376_ _12368_/X _12376_/B _12376_/C _12375_/X VGND VGND VPWR VPWR _12376_/X sky130_fd_sc_hd__or4_4
XANTENNA__22461__A3 _22459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20823__A _20802_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14115_ _14119_/A VGND VGND VPWR VPWR _14115_/X sky130_fd_sc_hd__buf_2
XFILLER_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15095_ _15158_/A VGND VGND VPWR VPWR _15144_/A sky130_fd_sc_hd__inv_2
X_19972_ _23141_/Q VGND VGND VPWR VPWR _21953_/B sky130_fd_sc_hd__inv_2
XFILLER_125_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14046_ _14046_/A VGND VGND VPWR VPWR _17197_/B sky130_fd_sc_hd__buf_2
X_18923_ _18919_/Y _18922_/X _18901_/X _18922_/X VGND VGND VPWR VPWR _23518_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18854_ _18854_/A VGND VGND VPWR VPWR _18854_/X sky130_fd_sc_hd__buf_2
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17805_ _17708_/X _17804_/X _23931_/Q _17767_/X VGND VGND VPWR VPWR _23931_/D sky130_fd_sc_hd__o22a_4
X_15997_ _24362_/Q VGND VGND VPWR VPWR _15997_/Y sky130_fd_sc_hd__inv_2
X_18785_ _18798_/A VGND VGND VPWR VPWR _18785_/X sky130_fd_sc_hd__buf_2
XFILLER_95_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15651__A2 _15647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21444__A2_N _20826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14948_ _24667_/Q VGND VGND VPWR VPWR _15177_/A sky130_fd_sc_hd__inv_2
X_17736_ _17782_/A _23589_/Q VGND VGND VPWR VPWR _17736_/X sky130_fd_sc_hd__or2_4
XFILLER_63_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_35_0_HCLK clkbuf_8_35_0_HCLK/A VGND VGND VPWR VPWR _23385_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18050__B1 _18049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15939__B1 _11548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14879_ _15004_/A _15003_/A _14879_/C _15003_/B VGND VGND VPWR VPWR _14879_/X sky130_fd_sc_hd__or4_4
X_17667_ _17662_/A _17662_/B _15807_/X VGND VGND VPWR VPWR _17667_/X sky130_fd_sc_hd__o21a_4
XFILLER_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_98_0_HCLK clkbuf_8_99_0_HCLK/A VGND VGND VPWR VPWR _24079_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_36_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24286__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19406_ _13217_/B VGND VGND VPWR VPWR _19406_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16618_ _16616_/Y _16570_/A _16617_/X _16570_/A VGND VGND VPWR VPWR _16618_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17598_ _17595_/C _17607_/B VGND VGND VPWR VPWR _17605_/B sky130_fd_sc_hd__or2_4
XFILLER_23_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24215__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22375__A1_N _20747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16549_ _16530_/A VGND VGND VPWR VPWR _16549_/X sky130_fd_sc_hd__buf_2
X_19337_ _19336_/Y _19334_/X _19221_/X _19334_/X VGND VGND VPWR VPWR _19337_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13900__A _13908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19268_ _21701_/D VGND VGND VPWR VPWR _19268_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18219_ _18207_/X _18263_/B VGND VGND VPWR VPWR _18219_/X sky130_fd_sc_hd__or2_4
XANTENNA__22437__B1 _20744_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19199_ _19198_/Y _19196_/X _19109_/X _19196_/X VGND VGND VPWR VPWR _23419_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14914__B2 _14913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21230_ _21387_/A _21227_/X _21230_/C VGND VGND VPWR VPWR _21230_/X sky130_fd_sc_hd__and3_4
XFILLER_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21161_ _18048_/X VGND VGND VPWR VPWR _21930_/A sky130_fd_sc_hd__buf_2
XANTENNA__20463__A2 _13506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23850__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25074__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20112_ _23087_/Q VGND VGND VPWR VPWR _20112_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21092_ _20861_/B _21092_/B VGND VGND VPWR VPWR _21275_/A sky130_fd_sc_hd__or2_4
XANTENNA__25003__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20043_ _23114_/Q VGND VGND VPWR VPWR _20043_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17616__B1 _16748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21412__A1 _22444_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24920_ _24923_/CLK _13696_/X HRESETn VGND VGND VPWR VPWR _24920_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21564__A _21564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24851_ _24851_/CLK _14118_/X HRESETn VGND VGND VPWR VPWR _14107_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_6_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19369__B1 _19232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15562__A _15561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22379__B _22379_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23802_ _23898_/CLK _18639_/X HRESETn VGND VGND VPWR VPWR _23802_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21176__B1 _21175_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24782_ _23618_/CLK _14318_/X HRESETn VGND VGND VPWR VPWR _20177_/C sky130_fd_sc_hd__dfrtp_4
X_21994_ _22646_/A VGND VGND VPWR VPWR _21994_/X sky130_fd_sc_hd__buf_2
XFILLER_22_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23733_ _24167_/CLK _20582_/Y HRESETn VGND VGND VPWR VPWR _13532_/A sky130_fd_sc_hd__dfrtp_4
X_20945_ _22084_/A _19733_/Y VGND VGND VPWR VPWR _20945_/X sky130_fd_sc_hd__or2_4
XPHY_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_6_0_HCLK clkbuf_5_6_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23664_ _23664_/CLK _20726_/X HRESETn VGND VGND VPWR VPWR _23666_/D sky130_fd_sc_hd__dfstp_4
X_20876_ _20875_/X VGND VGND VPWR VPWR _20876_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22395__A _22395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17489__A _17487_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22615_ _14737_/A _22574_/B VGND VGND VPWR VPWR _22619_/B sky130_fd_sc_hd__or2_4
XPHY_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16393__A _16043_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23595_ _23596_/CLK _18701_/X VGND VGND VPWR VPWR _23595_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16355__B1 _16093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22546_ _22546_/A VGND VGND VPWR VPWR _22546_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23938__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22477_ _22477_/A _22477_/B VGND VGND VPWR VPWR _22477_/Y sky130_fd_sc_hd__nor2_4
X_12230_ _12149_/Y _12229_/X VGND VGND VPWR VPWR _12230_/X sky130_fd_sc_hd__or2_4
X_24216_ _24213_/CLK _16410_/X HRESETn VGND VGND VPWR VPWR _24216_/Q sky130_fd_sc_hd__dfrtp_4
X_21428_ _21428_/A VGND VGND VPWR VPWR _21428_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21739__A _14206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25196_ _23986_/CLK _11617_/X HRESETn VGND VGND VPWR VPWR _11614_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12161_ _12131_/X _12140_/X _12161_/C _12161_/D VGND VGND VPWR VPWR _12162_/B sky130_fd_sc_hd__or4_4
XFILLER_29_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24147_ _24264_/CLK _16585_/X HRESETn VGND VGND VPWR VPWR _24147_/Q sky130_fd_sc_hd__dfrtp_4
X_21359_ _23104_/Q _14016_/A _23080_/Q _22042_/B VGND VGND VPWR VPWR _21359_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14133__A2 _14122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12092_ _12091_/Y _24545_/Q _12091_/Y _24545_/Q VGND VGND VPWR VPWR _12092_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24078_ _24412_/CLK _16897_/X HRESETn VGND VGND VPWR VPWR _16765_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_77_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15920_ _15920_/A _15919_/X VGND VGND VPWR VPWR _15921_/A sky130_fd_sc_hd__and2_4
X_23029_ _23028_/X VGND VGND VPWR VPWR _23029_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15851_ _24417_/Q VGND VGND VPWR VPWR _15851_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24797__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16568__A _16566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14802_ _15092_/A _24126_/Q _24687_/Q _14801_/Y VGND VGND VPWR VPWR _14802_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24726__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15782_ _15781_/X _15763_/X _16087_/A _22463_/A _15779_/X VGND VGND VPWR VPWR _24444_/D
+ sky130_fd_sc_hd__a32o_4
X_18570_ _16330_/Y _23835_/Q _16330_/Y _23835_/Q VGND VGND VPWR VPWR _18571_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_251_0_HCLK clkbuf_8_251_0_HCLK/A VGND VGND VPWR VPWR _24698_/CLK sky130_fd_sc_hd__clkbuf_1
X_12994_ _25010_/Q _12993_/Y VGND VGND VPWR VPWR _12994_/X sky130_fd_sc_hd__or2_4
XFILLER_18_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22174__A2_N _22637_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14733_ _24689_/Q _14732_/A _14844_/A _14732_/Y VGND VGND VPWR VPWR _14734_/D sky130_fd_sc_hd__o22a_4
X_17521_ _16733_/Y _17511_/X _17520_/X _17517_/B VGND VGND VPWR VPWR _17521_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22903__B2 _22657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11945_ _11944_/X VGND VGND VPWR VPWR _15422_/A sky130_fd_sc_hd__buf_2
XFILLER_55_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17452_ _17452_/A VGND VGND VPWR VPWR _17453_/A sky130_fd_sc_hd__inv_2
X_14664_ _14626_/A _14626_/B _14626_/A _14626_/B VGND VGND VPWR VPWR _14665_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11876_ _11871_/A _11873_/X _11874_/Y _11875_/Y VGND VGND VPWR VPWR _11876_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20818__A _20818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16403_ _16400_/Y _16396_/X _16243_/X _16402_/X VGND VGND VPWR VPWR _24219_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13615_ _13614_/X VGND VGND VPWR VPWR _21293_/B sky130_fd_sc_hd__buf_2
X_17383_ _17251_/Y _17382_/X _17336_/X VGND VGND VPWR VPWR _17383_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_60_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22667__B1 _14779_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14595_ _19144_/A _14589_/X _14594_/X VGND VGND VPWR VPWR _24734_/D sky130_fd_sc_hd__a21oi_4
X_16334_ HWDATA[21] VGND VGND VPWR VPWR _16334_/X sky130_fd_sc_hd__buf_2
X_19122_ _23446_/Q VGND VGND VPWR VPWR _19122_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13546_ _13546_/A VGND VGND VPWR VPWR _13546_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20101__A1_N _21931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12626__A2_N _24532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19053_ _13308_/B VGND VGND VPWR VPWR _19053_/Y sky130_fd_sc_hd__inv_2
X_16265_ _14929_/Y _16262_/X _16264_/X _16262_/X VGND VGND VPWR VPWR _24273_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23679__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13477_ _13475_/A _13480_/B _13476_/X VGND VGND VPWR VPWR _13478_/A sky130_fd_sc_hd__o21a_4
XANTENNA__22752__B _20807_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15216_ _15216_/A _15214_/Y _15226_/C VGND VGND VPWR VPWR _24656_/D sky130_fd_sc_hd__and3_4
X_18004_ _17999_/X _17990_/X _16558_/X _23910_/Q _17974_/X VGND VGND VPWR VPWR _23910_/D
+ sky130_fd_sc_hd__a32o_4
X_12428_ _12391_/Y _12425_/X _12419_/Y _12427_/X VGND VGND VPWR VPWR _12429_/A sky130_fd_sc_hd__a211o_4
XFILLER_126_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16196_ _16196_/A VGND VGND VPWR VPWR _16196_/X sky130_fd_sc_hd__buf_2
XFILLER_12_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20553__A _20552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15147_ _15144_/A VGND VGND VPWR VPWR _15147_/X sky130_fd_sc_hd__buf_2
XFILLER_127_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15647__A _15460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12359_ _25082_/Q VGND VGND VPWR VPWR _12360_/A sky130_fd_sc_hd__inv_2
XFILLER_47_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15078_ _15078_/A _15061_/B VGND VGND VPWR VPWR _15078_/Y sky130_fd_sc_hd__nand2_4
X_19955_ _19955_/A VGND VGND VPWR VPWR _19955_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12135__B2 _24568_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14029_ _14012_/Y _14026_/X _13663_/X _14028_/X VGND VGND VPWR VPWR _14029_/X sky130_fd_sc_hd__a2bb2o_4
X_18906_ _18899_/Y VGND VGND VPWR VPWR _18906_/X sky130_fd_sc_hd__buf_2
XFILLER_113_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19886_ _22075_/B _19885_/X _19815_/X _19885_/X VGND VGND VPWR VPWR _23174_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_61_0_HCLK clkbuf_6_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_61_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__21384__A _21224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18837_ _23548_/Q VGND VGND VPWR VPWR _18837_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24467__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18768_ _18768_/A VGND VGND VPWR VPWR _18768_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17719_ _17887_/A _17719_/B VGND VGND VPWR VPWR _17719_/X sky130_fd_sc_hd__or2_4
XFILLER_93_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18699_ _23595_/Q VGND VGND VPWR VPWR _18699_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20730_ _20729_/X VGND VGND VPWR VPWR _23662_/D sky130_fd_sc_hd__inv_2
XANTENNA__16585__B1 _16254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13399__B1 _13398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20661_ _23751_/Q _20660_/B _20660_/Y VGND VGND VPWR VPWR _20661_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_11_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14726__A _14726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22400_ _22226_/X _22399_/Y _14827_/Y _22228_/X VGND VGND VPWR VPWR _22400_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13630__A _16043_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20592_ _16534_/Y _20574_/X _20583_/X _20591_/Y VGND VGND VPWR VPWR _20592_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16337__B1 _16259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23380_ _23374_/CLK _23380_/D VGND VGND VPWR VPWR _13141_/B sky130_fd_sc_hd__dfxtp_4
X_22331_ _22495_/A _22321_/Y _22331_/C _22331_/D VGND VGND VPWR VPWR _22331_/X sky130_fd_sc_hd__or4_4
XFILLER_137_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24630__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25050_ _25050_/CLK _25050_/D HRESETn VGND VGND VPWR VPWR _12730_/A sky130_fd_sc_hd__dfrtp_4
X_22262_ _14047_/A _22256_/X _22258_/X _22262_/D VGND VGND VPWR VPWR _22262_/X sky130_fd_sc_hd__or4_4
XFILLER_105_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24001_ _25217_/CLK _17365_/X HRESETn VGND VGND VPWR VPWR _24001_/Q sky130_fd_sc_hd__dfrtp_4
X_21213_ _21238_/A VGND VGND VPWR VPWR _21214_/A sky130_fd_sc_hd__buf_2
XANTENNA__15557__A _15556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22193_ _16475_/A _22192_/X _22835_/A _25199_/Q _22858_/A VGND VGND VPWR VPWR _22193_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_117_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21144_ _21144_/A _21142_/X _21143_/X VGND VGND VPWR VPWR _21144_/X sky130_fd_sc_hd__and3_4
XFILLER_59_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21075_ _14302_/Y _12062_/X _24773_/Q _22018_/B VGND VGND VPWR VPWR _21075_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21397__B1 _21246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17065__A1 _17022_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20026_ _20026_/A VGND VGND VPWR VPWR _21326_/B sky130_fd_sc_hd__inv_2
XFILLER_115_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12412__C _12412_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24890__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24903_ _24902_/CLK _24903_/D HRESETn VGND VGND VPWR VPWR _24903_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24834_ _24851_/CLK _24834_/D HRESETn VGND VGND VPWR VPWR _12048_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18014__B1 _16617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24137__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11637__B1 _11636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24765_ _24851_/CLK _14398_/X HRESETn VGND VGND VPWR VPWR _14372_/A sky130_fd_sc_hd__dfrtp_4
X_21977_ _21050_/Y VGND VGND VPWR VPWR _22527_/B sky130_fd_sc_hd__buf_2
XPHY_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21904__A2_N _20818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11730_ _11729_/X VGND VGND VPWR VPWR _18065_/B sky130_fd_sc_hd__inv_2
XPHY_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23716_ _23716_/CLK _23716_/D HRESETn VGND VGND VPWR VPWR _20512_/A sky130_fd_sc_hd__dfrtp_4
X_20928_ _20900_/A VGND VGND VPWR VPWR _22488_/B sky130_fd_sc_hd__buf_2
XFILLER_70_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_81_0_HCLK clkbuf_8_81_0_HCLK/A VGND VGND VPWR VPWR _23624_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24696_ _24706_/CLK _15048_/Y HRESETn VGND VGND VPWR VPWR _14759_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20638__A _13537_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11661_ _24954_/Q VGND VGND VPWR VPWR _13591_/A sky130_fd_sc_hd__inv_2
XPHY_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23647_ _24783_/CLK _23647_/D HRESETn VGND VGND VPWR VPWR _20271_/A sky130_fd_sc_hd__dfstp_4
X_20859_ _18263_/A _20861_/B VGND VGND VPWR VPWR _20859_/X sky130_fd_sc_hd__and2_4
XPHY_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _24973_/Q VGND VGND VPWR VPWR _20883_/A sky130_fd_sc_hd__inv_2
XANTENNA__16591__A3 HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14380_ _13413_/Y _14380_/B VGND VGND VPWR VPWR _14380_/X sky130_fd_sc_hd__or2_4
XPHY_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11592_ _25202_/Q VGND VGND VPWR VPWR _11592_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21321__B1 _13334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23578_ _23563_/CLK _23578_/D VGND VGND VPWR VPWR _17864_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22853__A _22853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13331_ _20891_/A _13329_/Y _13330_/X _13329_/Y VGND VGND VPWR VPWR _13331_/X sky130_fd_sc_hd__a2bb2o_4
X_22529_ _17498_/A _22852_/A _13335_/X VGND VGND VPWR VPWR _22529_/X sky130_fd_sc_hd__a21o_4
XANTENNA__23772__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_HCLK clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16050_ _24353_/Q VGND VGND VPWR VPWR _16050_/Y sky130_fd_sc_hd__inv_2
X_13262_ _13166_/A _13262_/B VGND VGND VPWR VPWR _13263_/C sky130_fd_sc_hd__or2_4
XANTENNA__21469__A _21469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23701__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15001_ _15016_/A _14997_/B _15001_/C VGND VGND VPWR VPWR _15001_/X sky130_fd_sc_hd__or3_4
XFILLER_136_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12213_ _12186_/B _12184_/X _12185_/B VGND VGND VPWR VPWR _12213_/X sky130_fd_sc_hd__o21a_4
XFILLER_136_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13193_ _13057_/X _13192_/X _25000_/Q _13116_/X VGND VGND VPWR VPWR _25000_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21188__B _21187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25179_ _24847_/CLK _25179_/D HRESETn VGND VGND VPWR VPWR _11777_/A sky130_fd_sc_hd__dfrtp_4
X_12144_ _24573_/Q VGND VGND VPWR VPWR _12144_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24978__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16500__B1 _15484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17843__A3 _17842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19740_ _19740_/A VGND VGND VPWR VPWR _21925_/B sky130_fd_sc_hd__inv_2
XFILLER_2_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24907__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12075_ _12075_/A VGND VGND VPWR VPWR _12075_/Y sky130_fd_sc_hd__inv_2
X_16952_ _16778_/Y _16952_/B VGND VGND VPWR VPWR _16952_/Y sky130_fd_sc_hd__nand2_4
XFILLER_111_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21388__B1 _21231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15903_ _15902_/Y _15900_/X _15282_/X _15900_/X VGND VGND VPWR VPWR _15903_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14210__A1_N _20235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19671_ _21910_/B _19668_/X _19600_/X _19668_/X VGND VGND VPWR VPWR _23253_/D sky130_fd_sc_hd__a2bb2o_4
X_16883_ _16940_/A VGND VGND VPWR VPWR _16890_/A sky130_fd_sc_hd__buf_2
XFILLER_49_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16298__A _18263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14840__A1_N _24699_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24560__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18622_ _23642_/Q _18619_/X VGND VGND VPWR VPWR _18622_/X sky130_fd_sc_hd__or2_4
X_15834_ _15847_/A VGND VGND VPWR VPWR _15834_/X sky130_fd_sc_hd__buf_2
XFILLER_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21932__A _21342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18553_ _18422_/Y _18552_/X _18449_/X VGND VGND VPWR VPWR _18553_/Y sky130_fd_sc_hd__a21oi_4
X_12977_ _12774_/Y _12974_/X VGND VGND VPWR VPWR _12977_/X sky130_fd_sc_hd__or2_4
X_15765_ HWDATA[22] VGND VGND VPWR VPWR _15765_/X sky130_fd_sc_hd__buf_2
X_17504_ _17515_/D _17515_/B VGND VGND VPWR VPWR _17505_/D sky130_fd_sc_hd__or2_4
XFILLER_61_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11928_ _25160_/Q VGND VGND VPWR VPWR _11928_/Y sky130_fd_sc_hd__inv_2
X_14716_ _15096_/A VGND VGND VPWR VPWR _14716_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21651__B _21651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19402__A _19396_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15696_ _12316_/Y _15695_/X _13658_/X _15695_/X VGND VGND VPWR VPWR _15696_/X sky130_fd_sc_hd__a2bb2o_4
X_18484_ _18484_/A VGND VGND VPWR VPWR _18504_/A sky130_fd_sc_hd__buf_2
XFILLER_60_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16567__B1 _24156_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21560__B1 _21559_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14647_ _14620_/A VGND VGND VPWR VPWR _14647_/X sky130_fd_sc_hd__buf_2
X_17435_ _17264_/Y _17434_/X VGND VGND VPWR VPWR _17435_/X sky130_fd_sc_hd__or2_4
X_11859_ _25169_/Q VGND VGND VPWR VPWR _11859_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_109_0_HCLK clkbuf_7_54_0_HCLK/X VGND VGND VPWR VPWR _24013_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16582__A3 _15600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14578_ _14577_/X VGND VGND VPWR VPWR _17694_/A sky130_fd_sc_hd__buf_2
X_17366_ _17329_/A _17505_/C VGND VGND VPWR VPWR _17366_/X sky130_fd_sc_hd__and2_4
XANTENNA__16319__B1 _16246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19105_ _23452_/Q VGND VGND VPWR VPWR _19105_/Y sky130_fd_sc_hd__inv_2
X_13529_ _23730_/Q _13529_/B VGND VGND VPWR VPWR _13529_/X sky130_fd_sc_hd__or2_4
X_16317_ _16316_/Y _16314_/X _11536_/X _16314_/X VGND VGND VPWR VPWR _24250_/D sky130_fd_sc_hd__a2bb2o_4
X_17297_ _17297_/A _17296_/X VGND VGND VPWR VPWR _17586_/A sky130_fd_sc_hd__or2_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12066__A _16559_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16248_ _14901_/Y _16242_/X _16246_/X _16247_/X VGND VGND VPWR VPWR _24282_/D sky130_fd_sc_hd__a2bb2o_4
X_19036_ _19031_/Y _19035_/X _18901_/X _19035_/X VGND VGND VPWR VPWR _19036_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21379__A _21394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16179_ HWDATA[16] VGND VGND VPWR VPWR _16179_/X sky130_fd_sc_hd__buf_2
XFILLER_86_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24648__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19938_ _23153_/Q VGND VGND VPWR VPWR _19938_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22040__A1 _22146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19869_ _19876_/A VGND VGND VPWR VPWR _19869_/X sky130_fd_sc_hd__buf_2
XANTENNA__15824__B _16135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21900_ _21899_/X VGND VGND VPWR VPWR _21900_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13625__A _13624_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19992__B1 _17993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22880_ _24217_/Q _22806_/B VGND VGND VPWR VPWR _22880_/X sky130_fd_sc_hd__or2_4
XANTENNA__16001__A _24360_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22938__A _22997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24230__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21831_ _20946_/X _21831_/B VGND VGND VPWR VPWR _21831_/X sky130_fd_sc_hd__or2_4
XFILLER_71_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21842__A _12403_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16936__A _16936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19746__A2_N _19743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24550_ _24521_/CLK _24550_/D HRESETn VGND VGND VPWR VPWR _24550_/Q sky130_fd_sc_hd__dfrtp_4
X_21762_ _21234_/A VGND VGND VPWR VPWR _21762_/X sky130_fd_sc_hd__buf_2
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_68_0_HCLK clkbuf_6_34_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_68_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23501_ _23560_/CLK _23501_/D VGND VGND VPWR VPWR _13068_/B sky130_fd_sc_hd__dfxtp_4
X_20713_ _23624_/Q VGND VGND VPWR VPWR _20713_/Y sky130_fd_sc_hd__inv_2
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24481_ _24478_/CLK _15688_/X HRESETn VGND VGND VPWR VPWR _24481_/Q sky130_fd_sc_hd__dfrtp_4
X_21693_ _15430_/A _21692_/X _24929_/Q _15430_/A VGND VGND VPWR VPWR _21693_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12044__B1 _11985_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23432_ _23425_/CLK _19163_/X VGND VGND VPWR VPWR _23432_/Q sky130_fd_sc_hd__dfxtp_4
X_20644_ _20643_/Y _20644_/B VGND VGND VPWR VPWR _20644_/X sky130_fd_sc_hd__and2_4
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22649__A2_N _22643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23363_ _23350_/CLK _23363_/D VGND VGND VPWR VPWR _13175_/B sky130_fd_sc_hd__dfxtp_4
X_20575_ _23732_/Q VGND VGND VPWR VPWR _20575_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16671__A _16291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25102_ _25115_/CLK _12302_/Y HRESETn VGND VGND VPWR VPWR _25102_/Q sky130_fd_sc_hd__dfrtp_4
X_22314_ _16098_/Y _22314_/B VGND VGND VPWR VPWR _22314_/X sky130_fd_sc_hd__and2_4
XANTENNA__17486__B _21839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23294_ _23388_/CLK _23294_/D VGND VGND VPWR VPWR _23294_/Q sky130_fd_sc_hd__dfxtp_4
X_25033_ _25034_/CLK _25033_/D HRESETn VGND VGND VPWR VPWR _22921_/A sky130_fd_sc_hd__dfrtp_4
X_22245_ _22245_/A _22245_/B VGND VGND VPWR VPWR _22245_/X sky130_fd_sc_hd__and2_4
XFILLER_121_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22803__B1 _22351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22176_ _15463_/A VGND VGND VPWR VPWR _22857_/B sky130_fd_sc_hd__buf_2
XANTENNA__20921__A _22445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24389__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21127_ _21108_/X _21127_/B _21123_/Y _21127_/D VGND VGND VPWR VPWR _21127_/X sky130_fd_sc_hd__or4_4
XFILLER_120_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24318__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21058_ _22835_/A VGND VGND VPWR VPWR _21058_/X sky130_fd_sc_hd__buf_2
XFILLER_59_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12900_ _12899_/X VGND VGND VPWR VPWR _12900_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19983__B1 _15556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20009_ _20729_/B _23665_/Q VGND VGND VPWR VPWR _20010_/A sky130_fd_sc_hd__or2_4
X_13880_ _13852_/A _13880_/B _13880_/C VGND VGND VPWR VPWR _13881_/A sky130_fd_sc_hd__or3_4
XFILLER_98_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16797__B1 _24405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22848__A _24493_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12831_ _12964_/A _22365_/A _12964_/A _22365_/A VGND VGND VPWR VPWR _12835_/C sky130_fd_sc_hd__a2bb2o_4
X_24817_ _24788_/CLK _24817_/D HRESETn VGND VGND VPWR VPWR _24817_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16846__A _16846_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15550_ _19448_/A VGND VGND VPWR VPWR _15550_/X sky130_fd_sc_hd__buf_2
XFILLER_128_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12762_ _12651_/C _12735_/X VGND VGND VPWR VPWR _12762_/X sky130_fd_sc_hd__or2_4
X_24748_ _24748_/CLK _14518_/X HRESETn VGND VGND VPWR VPWR _21751_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14500_/Y _14480_/X _24749_/Q _14484_/X VGND VGND VPWR VPWR _14501_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16565__B _16235_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11698_/C _11704_/Y _11702_/X _11712_/X VGND VGND VPWR VPWR _25188_/D sky130_fd_sc_hd__o22a_4
XPHY_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _12101_/Y _15475_/X _11552_/X _15475_/X VGND VGND VPWR VPWR _15481_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23953__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12605_/A _12692_/Y VGND VGND VPWR VPWR _12693_/X sky130_fd_sc_hd__or2_4
X_24679_ _24681_/CLK _24679_/D HRESETn VGND VGND VPWR VPWR _24679_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25177__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _14432_/A _15449_/A VGND VGND VPWR VPWR _14432_/X sky130_fd_sc_hd__and2_4
X_17220_ _13613_/A _12061_/B _14013_/A VGND VGND VPWR VPWR _17220_/X sky130_fd_sc_hd__or3_4
XPHY_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11640_/Y _11521_/A _11643_/X _11521_/A VGND VGND VPWR VPWR _25190_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25106__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17151_ _17129_/A _17145_/B _17150_/Y VGND VGND VPWR VPWR _24034_/D sky130_fd_sc_hd__and3_4
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14363_ _14356_/X _14362_/Y sda_oen_o_S4 _14356_/X VGND VGND VPWR VPWR _24770_/D
+ sky130_fd_sc_hd__a2bb2o_4
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11575_ _11575_/A VGND VGND VPWR VPWR _11575_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16581__A _16581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16102_ _16102_/A VGND VGND VPWR VPWR _22267_/A sky130_fd_sc_hd__inv_2
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13314_ _13065_/X _13312_/X _13314_/C VGND VGND VPWR VPWR _13314_/X sky130_fd_sc_hd__and3_4
X_17082_ _17052_/A _17080_/X _17081_/X VGND VGND VPWR VPWR _24052_/D sky130_fd_sc_hd__and3_4
X_14294_ _14292_/Y _14288_/X _14236_/X _14293_/X VGND VGND VPWR VPWR _14294_/X sky130_fd_sc_hd__a2bb2o_4
X_16033_ _19144_/B _16033_/B VGND VGND VPWR VPWR _16033_/Y sky130_fd_sc_hd__nor2_4
X_13245_ _13309_/A _13245_/B VGND VGND VPWR VPWR _13245_/X sky130_fd_sc_hd__or2_4
XFILLER_108_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13176_ _13090_/X _13174_/X _13175_/X VGND VGND VPWR VPWR _13176_/X sky130_fd_sc_hd__and3_4
XFILLER_83_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11561__A2 _11535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12127_ _12127_/A VGND VGND VPWR VPWR _12127_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24741__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17984_ _17982_/X _15430_/X _11585_/A _22450_/A _17983_/X VGND VGND VPWR VPWR _23924_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_2_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24059__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19723_ _19723_/A VGND VGND VPWR VPWR _21459_/B sky130_fd_sc_hd__inv_2
X_12058_ _20695_/B _12057_/X SCLK_S3 _20695_/B VGND VGND VPWR VPWR _25136_/D sky130_fd_sc_hd__a2bb2o_4
X_16935_ _16935_/A _16938_/B VGND VGND VPWR VPWR _16935_/Y sky130_fd_sc_hd__nand2_4
XFILLER_46_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19654_ _19654_/A VGND VGND VPWR VPWR _19654_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16866_ _16866_/A _16866_/B VGND VGND VPWR VPWR _16866_/X sky130_fd_sc_hd__or2_4
XANTENNA__16788__B1 _24400_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18605_ _18604_/X VGND VGND VPWR VPWR _23812_/D sky130_fd_sc_hd__inv_2
X_15817_ _15720_/X _15815_/Y _15712_/X _15815_/Y VGND VGND VPWR VPWR _15817_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19585_ _19585_/A VGND VGND VPWR VPWR _21514_/B sky130_fd_sc_hd__inv_2
X_16797_ _15851_/Y _24081_/Q _24405_/Q _16834_/D VGND VGND VPWR VPWR _16804_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22477__B _22477_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15660__A _15664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18536_ _18536_/A _18536_/B VGND VGND VPWR VPWR _18536_/X sky130_fd_sc_hd__or2_4
XFILLER_34_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15748_ _16581_/A VGND VGND VPWR VPWR _15748_/X sky130_fd_sc_hd__buf_2
XANTENNA__16475__B _16475_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23694__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18467_ _18467_/A VGND VGND VPWR VPWR _23839_/D sky130_fd_sc_hd__inv_2
X_15679_ _12382_/Y _15677_/X _11563_/X _15677_/X VGND VGND VPWR VPWR _24487_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17418_ _17415_/A _17421_/B VGND VGND VPWR VPWR _17418_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__23623__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18398_ _16408_/Y _23839_/Q _24210_/Q _18488_/A VGND VGND VPWR VPWR _18401_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16960__B1 _16133_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17349_ _17349_/A _17349_/B VGND VGND VPWR VPWR _17358_/B sky130_fd_sc_hd__or2_4
XFILLER_105_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20360_ _17174_/X _20359_/Y _20349_/X VGND VGND VPWR VPWR _20360_/X sky130_fd_sc_hd__and3_4
XFILLER_31_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19019_ _21769_/B _19013_/X _15550_/X _19018_/X VGND VGND VPWR VPWR _23484_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24829__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20291_ _20291_/A VGND VGND VPWR VPWR _23632_/D sky130_fd_sc_hd__inv_2
X_22030_ _22030_/A _21106_/X VGND VGND VPWR VPWR _22030_/X sky130_fd_sc_hd__and2_4
XFILLER_115_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16743__A2_N _16685_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24482__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20811__A2 _20799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24411__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23981_ _25194_/CLK _17438_/X HRESETn VGND VGND VPWR VPWR _17318_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_130_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13373__A1_N _11890_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_31_0_HCLK clkbuf_5_30_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22932_ _20542_/B _22285_/X _23755_/Q _22531_/X VGND VGND VPWR VPWR _22932_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_110_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21572__A _24097_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22863_ _24216_/Q _23020_/B VGND VGND VPWR VPWR _22867_/B sky130_fd_sc_hd__or2_4
XANTENNA__16666__A _16643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15570__A _21292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24602_ _23744_/CLK _15360_/X HRESETn VGND VGND VPWR VPWR _15357_/A sky130_fd_sc_hd__dfrtp_4
X_21814_ _21810_/X _21813_/X _22105_/A VGND VGND VPWR VPWR _21814_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21291__B _20749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22794_ _22017_/X _22792_/X _21882_/X _22793_/X VGND VGND VPWR VPWR _22794_/X sky130_fd_sc_hd__o22a_4
XFILLER_25_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24533_ _24478_/CLK _24533_/D HRESETn VGND VGND VPWR VPWR _24533_/Q sky130_fd_sc_hd__dfrtp_4
X_21745_ _21564_/A _21723_/Y _21726_/X _21732_/Y _21744_/X VGND VGND VPWR VPWR _21745_/X
+ sky130_fd_sc_hd__a2111o_4
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14006__A1 _14004_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13090__A _11751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11603__A _25199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24464_ _23442_/CLK _24464_/D HRESETn VGND VGND VPWR VPWR _15716_/A sky130_fd_sc_hd__dfrtp_4
X_21676_ _21657_/A _21676_/B VGND VGND VPWR VPWR _21678_/B sky130_fd_sc_hd__or2_4
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23415_ _23419_/CLK _23415_/D VGND VGND VPWR VPWR _23415_/Q sky130_fd_sc_hd__dfxtp_4
X_20627_ _20627_/A VGND VGND VPWR VPWR _20627_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_155_0_HCLK clkbuf_7_77_0_HCLK/X VGND VGND VPWR VPWR _25005_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24395_ _24620_/CLK _15909_/X HRESETn VGND VGND VPWR VPWR _24395_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23346_ _23336_/CLK _23346_/D VGND VGND VPWR VPWR _13217_/B sky130_fd_sc_hd__dfxtp_4
X_20558_ _20558_/A VGND VGND VPWR VPWR _20558_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23277_ _23278_/CLK _19601_/X VGND VGND VPWR VPWR _19599_/A sky130_fd_sc_hd__dfxtp_4
X_20489_ _20484_/X _20487_/Y _24599_/Q _20488_/X VGND VGND VPWR VPWR _23710_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12434__A _12434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23663__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13030_ _13049_/A _13030_/B VGND VGND VPWR VPWR _13030_/X sky130_fd_sc_hd__or2_4
XFILLER_65_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25016_ _25034_/CLK _25016_/D HRESETn VGND VGND VPWR VPWR _22308_/A sky130_fd_sc_hd__dfrtp_4
X_22228_ _22228_/A VGND VGND VPWR VPWR _22228_/X sky130_fd_sc_hd__buf_2
XANTENNA__22252__A1 _15463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22252__B2 _15824_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20651__A _20651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18759__C _13461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22159_ _11961_/X VGND VGND VPWR VPWR _22952_/B sky130_fd_sc_hd__buf_2
XANTENNA__22526__A2_N _22523_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24152__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15464__B _15459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14981_ _15014_/A _14981_/B _14981_/C VGND VGND VPWR VPWR _14981_/X sky130_fd_sc_hd__and3_4
XANTENNA__19956__B1 _19381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15690__B1 _24480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16720_ _16720_/A VGND VGND VPWR VPWR _17489_/C sky130_fd_sc_hd__inv_2
X_13932_ _24895_/Q VGND VGND VPWR VPWR _13947_/A sky130_fd_sc_hd__inv_2
XFILLER_93_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13863_ _13863_/A _13897_/B _13862_/Y VGND VGND VPWR VPWR _14357_/C sky130_fd_sc_hd__or3_4
X_16651_ _16649_/Y _16650_/X _15497_/X _16650_/X VGND VGND VPWR VPWR _16651_/X sky130_fd_sc_hd__a2bb2o_4
X_12814_ _12812_/A _12813_/A _12812_/Y _12813_/Y VGND VGND VPWR VPWR _12821_/B sky130_fd_sc_hd__o22a_4
X_15602_ _12619_/Y _15593_/X _11558_/X _15593_/X VGND VGND VPWR VPWR _24524_/D sky130_fd_sc_hd__a2bb2o_4
X_19370_ _13028_/B VGND VGND VPWR VPWR _19370_/Y sky130_fd_sc_hd__inv_2
X_13794_ _13794_/A VGND VGND VPWR VPWR _13794_/Y sky130_fd_sc_hd__inv_2
X_16582_ _16581_/X _16573_/X _15600_/X _24148_/Q _16566_/X VGND VGND VPWR VPWR _16582_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_128_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18321_ _18321_/A VGND VGND VPWR VPWR _18322_/B sky130_fd_sc_hd__inv_2
X_12745_ _12649_/C _12747_/B _12744_/Y VGND VGND VPWR VPWR _25048_/D sky130_fd_sc_hd__o21a_4
X_15533_ _24541_/Q VGND VGND VPWR VPWR _19442_/A sky130_fd_sc_hd__buf_2
XFILLER_16_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_51_0_HCLK clkbuf_7_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_51_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15464_ _15463_/X _15459_/A VGND VGND VPWR VPWR _15464_/X sky130_fd_sc_hd__or2_4
X_18252_ _18242_/A _18250_/X _18251_/Y VGND VGND VPWR VPWR _23870_/D sky130_fd_sc_hd__o21a_4
XANTENNA__12008__B1 _11636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12676_ _12676_/A VGND VGND VPWR VPWR _12676_/Y sky130_fd_sc_hd__inv_2
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _14403_/A VGND VGND VPWR VPWR _14415_/X sky130_fd_sc_hd__buf_2
X_17203_ _17201_/Y _17198_/X _17202_/X _17198_/X VGND VGND VPWR VPWR _17203_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _11623_/Y _11621_/X _11626_/X _11621_/X VGND VGND VPWR VPWR _25194_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15395_ _15395_/A VGND VGND VPWR VPWR _15395_/Y sky130_fd_sc_hd__inv_2
X_18183_ _23867_/Q VGND VGND VPWR VPWR _18240_/C sky130_fd_sc_hd__inv_2
XANTENNA__16206__A1_N _16205_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ _24772_/Q _14325_/A _23077_/Q _14319_/X VGND VGND VPWR VPWR _14346_/X sky130_fd_sc_hd__o22a_4
X_17134_ _17134_/A _17154_/A VGND VGND VPWR VPWR _17134_/X sky130_fd_sc_hd__or2_4
XFILLER_50_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24993__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ HWDATA[22] VGND VGND VPWR VPWR _11558_/X sky130_fd_sc_hd__buf_2
XANTENNA__18695__B1 _17202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22491__A1 _23742_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22491__B2 _22170_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17065_ _17022_/B _17055_/B _17057_/X _17062_/B VGND VGND VPWR VPWR _17066_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24922__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14277_ _24795_/Q VGND VGND VPWR VPWR _14277_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21105__A2_N _11516_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16016_ _16014_/B _16014_/C VGND VGND VPWR VPWR _16016_/X sky130_fd_sc_hd__and2_4
X_13228_ _13122_/A _13226_/X _13227_/X VGND VGND VPWR VPWR _13228_/X sky130_fd_sc_hd__and3_4
XANTENNA__21735__A2_N _22439_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_14_0_HCLK_A clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15655__A _15655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13159_ _13075_/A VGND VGND VPWR VPWR _13159_/X sky130_fd_sc_hd__buf_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17967_ _17935_/A _18963_/A VGND VGND VPWR VPWR _17967_/X sky130_fd_sc_hd__or2_4
XFILLER_112_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15681__B1 _11566_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20006__B1 _19963_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19706_ _20972_/B _19701_/X _19641_/X _19688_/Y VGND VGND VPWR VPWR _23239_/D sky130_fd_sc_hd__a2bb2o_4
X_16918_ _16839_/B _16912_/X _16915_/B _16849_/X VGND VGND VPWR VPWR _16919_/A sky130_fd_sc_hd__a211o_4
X_17898_ _17898_/A _17898_/B _17898_/C VGND VGND VPWR VPWR _17898_/X sky130_fd_sc_hd__or3_4
XFILLER_22_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20557__B2 _20556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19637_ _21335_/B _19636_/X _19614_/X _19636_/X VGND VGND VPWR VPWR _23265_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16849_ _16858_/A VGND VGND VPWR VPWR _16849_/X sky130_fd_sc_hd__buf_2
XANTENNA__23875__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16486__A _16493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25099__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15390__A _16373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19568_ _21344_/B _19567_/X _11857_/X _19567_/X VGND VGND VPWR VPWR _23289_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23804__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22849__A3 _22839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25028__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18519_ _18504_/A _18519_/B _18519_/C VGND VGND VPWR VPWR _23826_/D sky130_fd_sc_hd__and3_4
XFILLER_94_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19499_ _19498_/Y _19494_/X _19455_/X _19494_/X VGND VGND VPWR VPWR _23314_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21530_ _21512_/X _21528_/X _21529_/X VGND VGND VPWR VPWR _21530_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_90_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22604__A1_N _21040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21461_ _21155_/A _21459_/X _21461_/C VGND VGND VPWR VPWR _21461_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_228_0_HCLK clkbuf_8_229_0_HCLK/A VGND VGND VPWR VPWR _24612_/CLK sky130_fd_sc_hd__clkbuf_1
X_23200_ _24008_/CLK _23200_/D VGND VGND VPWR VPWR _13269_/B sky130_fd_sc_hd__dfxtp_4
X_20412_ _15250_/X _20240_/X VGND VGND VPWR VPWR _23690_/D sky130_fd_sc_hd__and2_4
XANTENNA__18686__B1 _18685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24180_ _24180_/CLK _24180_/D HRESETn VGND VGND VPWR VPWR _24180_/Q sky130_fd_sc_hd__dfrtp_4
X_21392_ _21392_/A _21392_/B VGND VGND VPWR VPWR _21394_/B sky130_fd_sc_hd__or2_4
XFILLER_134_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12381__A2_N _21567_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24663__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23131_ _23128_/CLK _23131_/D VGND VGND VPWR VPWR _23131_/Q sky130_fd_sc_hd__dfxtp_4
X_20343_ _17187_/A VGND VGND VPWR VPWR _20343_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21567__A _21567_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23062_ _20740_/X VGND VGND VPWR VPWR IRQ[10] sky130_fd_sc_hd__buf_2
X_20274_ _23629_/Q _18624_/A VGND VGND VPWR VPWR _20274_/X sky130_fd_sc_hd__and2_4
XFILLER_103_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22013_ _20584_/Y _20749_/X _21867_/A _22012_/X VGND VGND VPWR VPWR _22013_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15565__A _19859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21286__B _21425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23964_ _24378_/CLK _23964_/D HRESETn VGND VGND VPWR VPWR _23964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22398__A _21246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20548__B2 _20465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22915_ _22914_/X VGND VGND VPWR VPWR _22915_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23895_ _23979_/CLK _23895_/D HRESETn VGND VGND VPWR VPWR _11757_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_112_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22846_ _22845_/X VGND VGND VPWR VPWR _22846_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12789__B2 _24455_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22777_ _15271_/A _22777_/B VGND VGND VPWR VPWR _22777_/Y sky130_fd_sc_hd__nor2_4
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _12536_/A _12536_/B VGND VGND VPWR VPWR _12537_/B sky130_fd_sc_hd__or2_4
Xclkbuf_6_38_0_HCLK clkbuf_6_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_76_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24516_ _24483_/CLK _24516_/D HRESETn VGND VGND VPWR VPWR _24516_/Q sky130_fd_sc_hd__dfrtp_4
X_21728_ _21728_/A _21425_/B VGND VGND VPWR VPWR _21728_/X sky130_fd_sc_hd__and2_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16843__B _16774_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12461_ _12415_/D _12424_/B _12415_/B VGND VGND VPWR VPWR _12461_/X sky130_fd_sc_hd__o21a_4
X_24447_ _24445_/CLK _24447_/D HRESETn VGND VGND VPWR VPWR _22595_/A sky130_fd_sc_hd__dfrtp_4
X_21659_ _21677_/A _21659_/B VGND VGND VPWR VPWR _21659_/X sky130_fd_sc_hd__or2_4
X_14200_ _14199_/B _14198_/X _14201_/A VGND VGND VPWR VPWR _14200_/X sky130_fd_sc_hd__a21o_4
X_15180_ _15165_/A _15177_/B _15180_/C VGND VGND VPWR VPWR _15180_/X sky130_fd_sc_hd__and3_4
X_12392_ _12391_/Y _22975_/A _12391_/Y _22975_/A VGND VGND VPWR VPWR _12396_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24378_ _24378_/CLK _15956_/X HRESETn VGND VGND VPWR VPWR _22598_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_126_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14131_ _13492_/X VGND VGND VPWR VPWR _14131_/X sky130_fd_sc_hd__buf_2
X_23329_ _23135_/CLK _23329_/D VGND VGND VPWR VPWR _19457_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_10_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24333__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14062_ _14062_/A VGND VGND VPWR VPWR _14062_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13013_ _13045_/A _13013_/B VGND VGND VPWR VPWR _13018_/B sky130_fd_sc_hd__or2_4
X_18870_ _18870_/A VGND VGND VPWR VPWR _18870_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17821_ _17821_/A _18721_/A VGND VGND VPWR VPWR _17821_/X sky130_fd_sc_hd__or2_4
XANTENNA__17652__A1 _21335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17690__A _14571_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11508__A _11507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17752_ _17898_/A _17746_/X _17752_/C VGND VGND VPWR VPWR _17764_/B sky130_fd_sc_hd__or3_4
X_14964_ _14964_/A VGND VGND VPWR VPWR _14964_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16703_ _22783_/A _22782_/A _15940_/Y _16702_/Y VGND VGND VPWR VPWR _16703_/X sky130_fd_sc_hd__o22a_4
X_13915_ _24898_/Q _13908_/X _13896_/X _24899_/Q _13911_/X VGND VGND VPWR VPWR _13915_/X
+ sky130_fd_sc_hd__a32o_4
X_17683_ _17676_/X _17681_/X _17682_/X VGND VGND VPWR VPWR _17683_/X sky130_fd_sc_hd__and3_4
X_14895_ _14895_/A VGND VGND VPWR VPWR _15179_/A sky130_fd_sc_hd__buf_2
XANTENNA__25192__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19422_ _19420_/Y _19418_/X _19421_/X _19418_/X VGND VGND VPWR VPWR _19422_/X sky130_fd_sc_hd__a2bb2o_4
X_16634_ _16624_/X _16625_/X HWDATA[26] _22857_/A _16622_/X VGND VGND VPWR VPWR _24119_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_74_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13846_ _13808_/X _13810_/X _13845_/A _13811_/B VGND VGND VPWR VPWR _13846_/X sky130_fd_sc_hd__or4_4
XANTENNA__11543__A2_N _11521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25121__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19353_ _19352_/Y _19350_/X _19308_/X _19350_/X VGND VGND VPWR VPWR _23365_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21940__A _21229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13777_ _13797_/A _14073_/B _13777_/C _13777_/D VGND VGND VPWR VPWR _13777_/X sky130_fd_sc_hd__or4_4
X_16565_ _22228_/A _16235_/B VGND VGND VPWR VPWR _16566_/A sky130_fd_sc_hd__or2_4
X_18304_ _18316_/A _18303_/X VGND VGND VPWR VPWR _18304_/X sky130_fd_sc_hd__or2_4
XFILLER_43_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15516_ _12104_/Y _15514_/X _15386_/X _15514_/X VGND VGND VPWR VPWR _15516_/X sky130_fd_sc_hd__a2bb2o_4
X_12728_ _12728_/A _12728_/B VGND VGND VPWR VPWR _12728_/X sky130_fd_sc_hd__or2_4
X_19284_ _19283_/Y VGND VGND VPWR VPWR _19284_/X sky130_fd_sc_hd__buf_2
XFILLER_31_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16496_ _16495_/Y _16493_/X _16251_/X _16493_/X VGND VGND VPWR VPWR _16496_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20556__A _20647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18235_ _18222_/B _18232_/X VGND VGND VPWR VPWR _18235_/X sky130_fd_sc_hd__or2_4
X_12659_ _25068_/Q _12658_/Y VGND VGND VPWR VPWR _12659_/X sky130_fd_sc_hd__or2_4
X_15447_ _14432_/X _15449_/B VGND VGND VPWR VPWR _15447_/X sky130_fd_sc_hd__and2_4
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18166_ _16080_/A _18278_/A _21716_/A _18322_/A VGND VGND VPWR VPWR _18172_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15378_ _24594_/Q VGND VGND VPWR VPWR _22278_/A sky130_fd_sc_hd__inv_2
XFILLER_106_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17117_ _17116_/X VGND VGND VPWR VPWR _17117_/Y sky130_fd_sc_hd__inv_2
X_14329_ _14329_/A _14329_/B VGND VGND VPWR VPWR _14329_/X sky130_fd_sc_hd__or2_4
X_18097_ _18104_/A _18104_/B _18096_/Y VGND VGND VPWR VPWR _18097_/X sky130_fd_sc_hd__a21o_4
XANTENNA__24074__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_58_0_HCLK clkbuf_8_59_0_HCLK/A VGND VGND VPWR VPWR _23992_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22216__A1 _20918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17048_ _17021_/Y _17055_/A _17067_/A _17054_/A VGND VGND VPWR VPWR _17048_/X sky130_fd_sc_hd__or4_4
XANTENNA__23809__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24003__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19093__B1 _18959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21975__B1 _12075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18999_ _21655_/B _18996_/X _15554_/X _18996_/X VGND VGND VPWR VPWR _23491_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25209__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16928__B _16927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20961_ _20961_/A _19684_/Y VGND VGND VPWR VPWR _20962_/C sky130_fd_sc_hd__or2_4
XANTENNA__22011__A _22011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15406__B1 _15291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22700_ _24488_/Q _22757_/B VGND VGND VPWR VPWR _22700_/X sky130_fd_sc_hd__or2_4
XFILLER_26_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23680_ _23680_/CLK _20401_/Y HRESETn VGND VGND VPWR VPWR _17186_/A sky130_fd_sc_hd__dfrtp_4
X_20892_ _22018_/B VGND VGND VPWR VPWR _20892_/X sky130_fd_sc_hd__buf_2
X_22631_ _22702_/A _22631_/B VGND VGND VPWR VPWR _22631_/X sky130_fd_sc_hd__and2_4
XANTENNA__22152__B1 _15430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22562_ _22677_/A _22562_/B _22562_/C VGND VGND VPWR VPWR _22572_/A sky130_fd_sc_hd__and3_4
XANTENNA__20466__A _20465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24301_ _24031_/CLK _24301_/D HRESETn VGND VGND VPWR VPWR _16188_/A sky130_fd_sc_hd__dfrtp_4
X_21513_ _21385_/A _21513_/B VGND VGND VPWR VPWR _21513_/X sky130_fd_sc_hd__or2_4
XFILLER_10_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24844__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22493_ _22175_/A _22491_/Y _22349_/B _22492_/X VGND VGND VPWR VPWR _22493_/X sky130_fd_sc_hd__o22a_4
XFILLER_22_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24232_ _23840_/CLK _16362_/X HRESETn VGND VGND VPWR VPWR _24232_/Q sky130_fd_sc_hd__dfrtp_4
X_21444_ _20332_/A _20826_/X _24811_/Q _21113_/C VGND VGND VPWR VPWR _21444_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21258__A2 _21255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22681__A _22681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24163_ _24162_/CLK _24163_/D HRESETn VGND VGND VPWR VPWR _16541_/A sky130_fd_sc_hd__dfrtp_4
X_21375_ _21211_/A _21375_/B VGND VGND VPWR VPWR _21375_/X sky130_fd_sc_hd__or2_4
X_23114_ _23292_/CLK _23114_/D VGND VGND VPWR VPWR _23114_/Q sky130_fd_sc_hd__dfxtp_4
X_20326_ _18619_/A _18619_/B _18620_/Y VGND VGND VPWR VPWR _20326_/Y sky130_fd_sc_hd__a21oi_4
X_24094_ _24094_/CLK _24094_/D HRESETn VGND VGND VPWR VPWR _14754_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19990__A _19989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23045_ VGND VGND VPWR VPWR _23045_/HI IRQ[13] sky130_fd_sc_hd__conb_1
X_20257_ _20225_/X _20257_/B _20244_/X _20257_/D VGND VGND VPWR VPWR _20257_/X sky130_fd_sc_hd__or4_4
XFILLER_135_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20769__A1 _20757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23797__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20188_ _20188_/A _13890_/A VGND VGND VPWR VPWR _20189_/B sky130_fd_sc_hd__and2_4
XFILLER_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23726__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24996_ _25002_/CLK _24996_/D HRESETn VGND VGND VPWR VPWR _24996_/Q sky130_fd_sc_hd__dfrtp_4
X_11961_ _13333_/A VGND VGND VPWR VPWR _11961_/X sky130_fd_sc_hd__buf_2
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23947_ _23972_/CLK _23947_/D HRESETn VGND VGND VPWR VPWR _23947_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13700_ _24918_/Q _13687_/X _24917_/Q _13689_/X VGND VGND VPWR VPWR _13700_/X sky130_fd_sc_hd__o22a_4
XFILLER_84_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22930__A2 _16134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14680_ _14609_/A VGND VGND VPWR VPWR _14680_/Y sky130_fd_sc_hd__inv_2
X_11892_ _11890_/A _11891_/A _11890_/Y _11891_/Y VGND VGND VPWR VPWR _11902_/A sky130_fd_sc_hd__o22a_4
XFILLER_45_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23878_ _25141_/CLK _18129_/X HRESETn VGND VGND VPWR VPWR _20886_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_72_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22856__A _22982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13631_ _13630_/X VGND VGND VPWR VPWR _13631_/X sky130_fd_sc_hd__buf_2
XFILLER_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22829_ _20527_/Y _22610_/X _23752_/Q _22657_/X VGND VGND VPWR VPWR _22829_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22143__B1 _22314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13562_ _13585_/A _13562_/B VGND VGND VPWR VPWR _13562_/X sky130_fd_sc_hd__or2_4
X_16350_ _16349_/Y _16347_/X _16087_/X _16347_/X VGND VGND VPWR VPWR _24237_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22694__A1 _24243_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12513_ _12512_/X VGND VGND VPWR VPWR _25080_/D sky130_fd_sc_hd__inv_2
X_15301_ _15300_/Y VGND VGND VPWR VPWR _15301_/X sky130_fd_sc_hd__buf_2
X_16281_ _14923_/Y _16278_/X _15978_/X _16278_/X VGND VGND VPWR VPWR _16281_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24585__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13493_ _24965_/Q _13388_/X _13488_/X VGND VGND VPWR VPWR _13521_/A sky130_fd_sc_hd__a21o_4
X_18020_ _19531_/A VGND VGND VPWR VPWR _18020_/X sky130_fd_sc_hd__buf_2
X_12444_ _12444_/A _12444_/B _12443_/X VGND VGND VPWR VPWR _12444_/X sky130_fd_sc_hd__or3_4
X_15232_ _14903_/Y _15123_/X _15126_/X _15230_/B VGND VGND VPWR VPWR _15232_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22446__A1 _24269_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24514__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_211_0_HCLK clkbuf_8_211_0_HCLK/A VGND VGND VPWR VPWR _24197_/CLK sky130_fd_sc_hd__clkbuf_1
X_15163_ _24671_/Q _15163_/B VGND VGND VPWR VPWR _15165_/B sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_3_0_0_HCLK_A clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12375_ _12489_/A _24482_/Q _12489_/A _24482_/Q VGND VGND VPWR VPWR _12375_/X sky130_fd_sc_hd__a2bb2o_4
X_14114_ _14111_/C _14110_/X VGND VGND VPWR VPWR _14119_/A sky130_fd_sc_hd__or2_4
X_15094_ _15094_/A VGND VGND VPWR VPWR _15158_/A sky130_fd_sc_hd__buf_2
X_19971_ _19967_/Y _19970_/X _19442_/A _19970_/X VGND VGND VPWR VPWR _19971_/X sky130_fd_sc_hd__a2bb2o_4
X_14045_ _14045_/A VGND VGND VPWR VPWR _14045_/Y sky130_fd_sc_hd__inv_2
X_18922_ _18935_/A VGND VGND VPWR VPWR _18922_/X sky130_fd_sc_hd__buf_2
XFILLER_106_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18853_ _18852_/X VGND VGND VPWR VPWR _18854_/A sky130_fd_sc_hd__inv_2
XANTENNA__21421__A2 _21553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17804_ _15730_/X _17785_/X _17803_/X _23932_/Q _17765_/X VGND VGND VPWR VPWR _17804_/X
+ sky130_fd_sc_hd__o32a_4
X_18784_ _18784_/A VGND VGND VPWR VPWR _18798_/A sky130_fd_sc_hd__inv_2
XFILLER_67_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15996_ _15995_/Y _15993_/X _15282_/X _15993_/X VGND VGND VPWR VPWR _15996_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17735_ _17721_/A VGND VGND VPWR VPWR _17782_/A sky130_fd_sc_hd__buf_2
XANTENNA__15651__A3 _15635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14947_ _14946_/Y _24278_/Q _14946_/Y _24278_/Q VGND VGND VPWR VPWR _14947_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21185__B2 _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17666_ _17665_/X VGND VGND VPWR VPWR _17666_/Y sky130_fd_sc_hd__inv_2
X_14878_ _14878_/A _14877_/X VGND VGND VPWR VPWR _15003_/B sky130_fd_sc_hd__or2_4
XANTENNA__20932__A1 _20550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19405_ _19404_/Y _19402_/X _19381_/X _19402_/X VGND VGND VPWR VPWR _23347_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16617_ _16216_/A VGND VGND VPWR VPWR _16617_/X sky130_fd_sc_hd__buf_2
XFILLER_1_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13829_ _13808_/A _13810_/A _24903_/Q _24902_/Q VGND VGND VPWR VPWR _13829_/X sky130_fd_sc_hd__or4_4
X_17597_ _17597_/A VGND VGND VPWR VPWR _17597_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19336_ _23371_/Q VGND VGND VPWR VPWR _19336_/Y sky130_fd_sc_hd__inv_2
X_16548_ _16548_/A VGND VGND VPWR VPWR _16548_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18889__B1 _18795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20286__A _13934_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_21_0_HCLK clkbuf_6_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19267_ _19265_/Y _19261_/X _19152_/X _19266_/X VGND VGND VPWR VPWR _23396_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16479_ _16479_/A VGND VGND VPWR VPWR _16530_/A sky130_fd_sc_hd__buf_2
X_18218_ _18295_/A _18218_/B _18218_/C VGND VGND VPWR VPWR _18263_/B sky130_fd_sc_hd__or3_4
XANTENNA__24255__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19198_ _23419_/Q VGND VGND VPWR VPWR _19198_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22988__A2 _22311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18149_ _24332_/Q _23853_/Q _16107_/Y _18210_/B VGND VGND VPWR VPWR _18149_/X sky130_fd_sc_hd__o22a_4
XFILLER_85_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21160_ _21346_/A _21160_/B _21160_/C VGND VGND VPWR VPWR _21160_/X sky130_fd_sc_hd__and3_4
XANTENNA__22006__A _22006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20111_ _20109_/Y _20110_/X _19614_/A _20110_/X VGND VGND VPWR VPWR _23088_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13628__A _22018_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21091_ _21072_/X _21078_/Y _21080_/Y _21090_/X VGND VGND VPWR VPWR _21091_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17616__A1 _17487_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20042_ _21831_/B _20036_/X _19717_/X _20041_/X VGND VGND VPWR VPWR _20042_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21845__A _24472_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23890__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15627__B1 _15390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24850_ _24968_/CLK _24850_/D HRESETn VGND VGND VPWR VPWR _14108_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_6_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21551__A2_N _23025_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25043__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19369__B2 _19349_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23801_ _24841_/CLK MSI_S3 HRESETn VGND VGND VPWR VPWR _23801_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24781_ _23618_/CLK _14323_/X HRESETn VGND VGND VPWR VPWR _20177_/A sky130_fd_sc_hd__dfrtp_4
X_21993_ _24366_/Q _22524_/B VGND VGND VPWR VPWR _21993_/X sky130_fd_sc_hd__or2_4
XANTENNA__16667__A1_N _14699_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23732_ _24162_/CLK _20578_/Y HRESETn VGND VGND VPWR VPWR _23732_/Q sky130_fd_sc_hd__dfrtp_4
X_20944_ _20971_/A VGND VGND VPWR VPWR _22084_/A sky130_fd_sc_hd__buf_2
XFILLER_82_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20923__A1 _21179_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11664__B2 _23913_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20923__B2 _12062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_103_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_207_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ _23664_/CLK _20724_/X HRESETn VGND VGND VPWR VPWR _23665_/D sky130_fd_sc_hd__dfstp_4
X_20875_ _20869_/X _20871_/X _20873_/X _20875_/D VGND VGND VPWR VPWR _20875_/X sky130_fd_sc_hd__or4_4
XPHY_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22614_ _22614_/A _22614_/B _22661_/C _22613_/X VGND VGND VPWR VPWR HRDATA[18] sky130_fd_sc_hd__or4_4
XANTENNA__22676__A1 _24415_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17489__B _17615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23594_ _23596_/CLK _18703_/X VGND VGND VPWR VPWR _18702_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16393__B _23763_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22545_ _21529_/X _22543_/X _13362_/A _22544_/X VGND VGND VPWR VPWR _22546_/A sky130_fd_sc_hd__o22a_4
XANTENNA__11611__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22476_ _21246_/X _22473_/X _22474_/X _22476_/D VGND VGND VPWR VPWR _22476_/X sky130_fd_sc_hd__or4_4
XANTENNA__12304__A1_N _12508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24215_ _24213_/CLK _24215_/D HRESETn VGND VGND VPWR VPWR _24215_/Q sky130_fd_sc_hd__dfrtp_4
X_21427_ _13335_/X _21423_/X _22407_/A _21426_/X VGND VGND VPWR VPWR _21428_/A sky130_fd_sc_hd__o22a_4
X_25195_ _25194_/CLK _11622_/X HRESETn VGND VGND VPWR VPWR _25195_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21739__B _21082_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12160_ _12153_/X _12160_/B _12160_/C _12159_/X VGND VGND VPWR VPWR _12161_/D sky130_fd_sc_hd__or4_4
X_24146_ _24145_/CLK _16586_/X HRESETn VGND VGND VPWR VPWR _24146_/Q sky130_fd_sc_hd__dfrtp_4
X_21358_ _15642_/X VGND VGND VPWR VPWR _22042_/B sky130_fd_sc_hd__buf_2
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14945__A2_N _22399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23978__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_41_0_HCLK clkbuf_7_20_0_HCLK/X VGND VGND VPWR VPWR _23511_/CLK sky130_fd_sc_hd__clkbuf_1
X_20309_ _20309_/A VGND VGND VPWR VPWR _23636_/D sky130_fd_sc_hd__inv_2
X_12091_ _25102_/Q VGND VGND VPWR VPWR _12091_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23907__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24077_ _24079_/CLK _16901_/X HRESETn VGND VGND VPWR VPWR _16780_/A sky130_fd_sc_hd__dfrtp_4
X_21289_ _21288_/X VGND VGND VPWR VPWR _21324_/B sky130_fd_sc_hd__inv_2
XFILLER_1_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23028_ _22429_/B _23024_/Y _22584_/A _23027_/X VGND VGND VPWR VPWR _23028_/X sky130_fd_sc_hd__o22a_4
XFILLER_131_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15618__B1 _24514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16849__A _16858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15753__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15850_ _15849_/Y _15847_/X _11555_/X _15847_/X VGND VGND VPWR VPWR _15850_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18173__A1_N _22401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14801_ _24130_/Q VGND VGND VPWR VPWR _14801_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21061__A1_N _21040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15781_ _16581_/A VGND VGND VPWR VPWR _15781_/X sky130_fd_sc_hd__buf_2
X_12993_ _12973_/B VGND VGND VPWR VPWR _12993_/Y sky130_fd_sc_hd__inv_2
X_24979_ _25141_/CLK _13378_/X HRESETn VGND VGND VPWR VPWR _13376_/A sky130_fd_sc_hd__dfrtp_4
X_17520_ _16747_/Y VGND VGND VPWR VPWR _17520_/X sky130_fd_sc_hd__buf_2
XFILLER_79_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13273__A _13136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14732_ _14732_/A VGND VGND VPWR VPWR _14732_/Y sky130_fd_sc_hd__inv_2
X_11944_ _22477_/B VGND VGND VPWR VPWR _11944_/X sky130_fd_sc_hd__buf_2
XFILLER_44_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17451_ _23976_/Q VGND VGND VPWR VPWR _17451_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24766__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11875_ _11871_/A _11871_/B _11868_/Y VGND VGND VPWR VPWR _11875_/Y sky130_fd_sc_hd__a21oi_4
X_14663_ _14655_/X _14662_/Y _24723_/Q _14655_/X VGND VGND VPWR VPWR _14663_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18188__A1_N _16054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16402_ _16426_/A VGND VGND VPWR VPWR _16402_/X sky130_fd_sc_hd__buf_2
X_13614_ _13614_/A VGND VGND VPWR VPWR _13614_/X sky130_fd_sc_hd__buf_2
X_17382_ _17266_/Y _17270_/Y _17382_/C _17382_/D VGND VGND VPWR VPWR _17382_/X sky130_fd_sc_hd__or4_4
X_14594_ _18719_/A VGND VGND VPWR VPWR _14594_/X sky130_fd_sc_hd__buf_2
X_19121_ _19119_/Y _19114_/X _19120_/X _19114_/A VGND VGND VPWR VPWR _19121_/X sky130_fd_sc_hd__a2bb2o_4
X_16333_ _16339_/A VGND VGND VPWR VPWR _16333_/X sky130_fd_sc_hd__buf_2
X_13545_ _23067_/Q _20554_/B VGND VGND VPWR VPWR _13545_/X sky130_fd_sc_hd__and2_4
XANTENNA__12080__B2 _24570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19052_ _19051_/Y _19049_/X _18938_/X _19049_/X VGND VGND VPWR VPWR _23472_/D sky130_fd_sc_hd__a2bb2o_4
X_13476_ _13403_/Y _13480_/A _13480_/A _13475_/Y VGND VGND VPWR VPWR _13476_/X sky130_fd_sc_hd__o22a_4
X_16264_ HWDATA[18] VGND VGND VPWR VPWR _16264_/X sky130_fd_sc_hd__buf_2
X_18003_ _11677_/Y _17987_/A _16617_/X _17987_/A VGND VGND VPWR VPWR _23911_/D sky130_fd_sc_hd__a2bb2o_4
X_12427_ _12442_/A VGND VGND VPWR VPWR _12427_/X sky130_fd_sc_hd__buf_2
X_15215_ _15158_/A VGND VGND VPWR VPWR _15226_/C sky130_fd_sc_hd__buf_2
XFILLER_138_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16195_ _16195_/A VGND VGND VPWR VPWR _16195_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12358_ _21104_/A _12356_/Y _25075_/Q _12357_/Y VGND VGND VPWR VPWR _12365_/B sky130_fd_sc_hd__a2bb2o_4
X_15146_ _15138_/B _15154_/B VGND VGND VPWR VPWR _15146_/X sky130_fd_sc_hd__or2_4
XANTENNA__11591__B1 _11590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15077_ _15057_/X _15071_/B _15077_/C VGND VGND VPWR VPWR _24689_/D sky130_fd_sc_hd__and3_4
X_19954_ _19952_/Y _19948_/X _19424_/X _19953_/X VGND VGND VPWR VPWR _19954_/X sky130_fd_sc_hd__a2bb2o_4
X_12289_ _12180_/B _12265_/X _12287_/B _12203_/X VGND VGND VPWR VPWR _12290_/A sky130_fd_sc_hd__a211o_4
XANTENNA__23648__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14028_ _14027_/X VGND VGND VPWR VPWR _14028_/X sky130_fd_sc_hd__buf_2
X_18905_ _23524_/Q VGND VGND VPWR VPWR _18905_/Y sky130_fd_sc_hd__inv_2
X_19885_ _19897_/A VGND VGND VPWR VPWR _19885_/X sky130_fd_sc_hd__buf_2
XFILLER_122_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15609__B1 _11570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18836_ _21947_/B _18833_/X _15545_/X _18833_/X VGND VGND VPWR VPWR _18836_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18767_ _18766_/Y _18762_/X _18740_/X _18762_/X VGND VGND VPWR VPWR _18767_/X sky130_fd_sc_hd__a2bb2o_4
X_15979_ _15987_/A VGND VGND VPWR VPWR _15979_/X sky130_fd_sc_hd__buf_2
XFILLER_3_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14832__B2 _14831_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17718_ _17727_/A VGND VGND VPWR VPWR _17887_/A sky130_fd_sc_hd__buf_2
XFILLER_23_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18698_ _18696_/Y _18692_/X _17205_/X _18697_/X VGND VGND VPWR VPWR _18698_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20905__A1 _21716_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20905__B2 _22859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17649_ _21144_/A _17648_/X _17626_/X _17630_/B VGND VGND VPWR VPWR _23939_/D sky130_fd_sc_hd__a22oi_4
XFILLER_51_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20728__B _23665_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24436__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20660_ _23751_/Q _20660_/B VGND VGND VPWR VPWR _20660_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__22658__B2 _22657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19319_ _19304_/Y VGND VGND VPWR VPWR _19319_/X sky130_fd_sc_hd__buf_2
XANTENNA__13630__B _23763_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20591_ _20590_/A _20590_/B _20590_/Y VGND VGND VPWR VPWR _20591_/Y sky130_fd_sc_hd__a21oi_4
X_22330_ _22330_/A VGND VGND VPWR VPWR _22331_/D sky130_fd_sc_hd__inv_2
XFILLER_30_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20744__A _20800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14899__B2 _24281_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22261_ _12406_/Y _22259_/X _16966_/A _22260_/X VGND VGND VPWR VPWR _22262_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19287__B1 _11839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24000_ _25217_/CLK _24000_/D HRESETn VGND VGND VPWR VPWR _24000_/Q sky130_fd_sc_hd__dfrtp_4
X_21212_ _21376_/A _21209_/X _21212_/C VGND VGND VPWR VPWR _21212_/X sky130_fd_sc_hd__and3_4
XANTENNA__21094__B1 _16616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22192_ _22192_/A _22439_/B VGND VGND VPWR VPWR _22192_/X sky130_fd_sc_hd__or2_4
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15848__B1 _15761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11582__B1 _11581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_0_0_HCLK clkbuf_8_1_0_HCLK/A VGND VGND VPWR VPWR _23100_/CLK sky130_fd_sc_hd__clkbuf_1
X_21143_ _21336_/A _19682_/Y VGND VGND VPWR VPWR _21143_/X sky130_fd_sc_hd__or2_4
XANTENNA__13358__A _13357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19039__B1 _19038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_28_0_HCLK clkbuf_6_14_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_28_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21074_ _14004_/Y _13333_/A _24801_/Q _11529_/A VGND VGND VPWR VPWR _21074_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20025_ _21460_/B _20020_/X _19724_/X _20020_/X VGND VGND VPWR VPWR _23121_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15573__A _22223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24902_ _24902_/CLK _13912_/X HRESETn VGND VGND VPWR VPWR _24902_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17491__C _16685_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16273__B1 _24269_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15615__A3 _15499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24833_ _24851_/CLK _24833_/D HRESETn VGND VGND VPWR VPWR _12048_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_73_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18884__A _18876_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13093__A _13169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21976_ _22702_/A _21975_/X VGND VGND VPWR VPWR _21976_/X sky130_fd_sc_hd__and2_4
XFILLER_55_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24764_ _24968_/CLK _24764_/D HRESETn VGND VGND VPWR VPWR _13416_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_54_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20919__A _20919_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20927_ _20926_/X VGND VGND VPWR VPWR _20927_/X sky130_fd_sc_hd__buf_2
XFILLER_14_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23715_ _23716_/CLK _23715_/D HRESETn VGND VGND VPWR VPWR _20513_/B sky130_fd_sc_hd__dfrtp_4
XPHY_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24695_ _24706_/CLK _15054_/X HRESETn VGND VGND VPWR VPWR _24695_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24177__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11660_ _11652_/X _11654_/X _11656_/X _11659_/X VGND VGND VPWR VPWR _11660_/X sky130_fd_sc_hd__or4_4
XPHY_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20858_ _24222_/Q _21273_/A _22153_/B _20857_/X VGND VGND VPWR VPWR _20858_/X sky130_fd_sc_hd__a211o_4
XPHY_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23646_ _23641_/CLK _23645_/Q HRESETn VGND VGND VPWR VPWR _23646_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_39_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24106__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13540__B _13539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11591_ _11587_/Y _11588_/X _11590_/X _11588_/X VGND VGND VPWR VPWR _25203_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17012__B _17007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23577_ _23568_/CLK _23577_/D VGND VGND VPWR VPWR _23577_/Q sky130_fd_sc_hd__dfxtp_4
X_20789_ _15407_/A VGND VGND VPWR VPWR _20826_/A sky130_fd_sc_hd__buf_2
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21321__B2 _21320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ _11643_/A VGND VGND VPWR VPWR _13330_/X sky130_fd_sc_hd__buf_2
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22528_ _12474_/C _22259_/A _17041_/A _22121_/X VGND VGND VPWR VPWR _22528_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ _13261_/A _23496_/Q VGND VGND VPWR VPWR _13261_/X sky130_fd_sc_hd__or2_4
XFILLER_109_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15748__A _16581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23030__A _22997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22459_ _22646_/A VGND VGND VPWR VPWR _22459_/X sky130_fd_sc_hd__buf_2
XANTENNA__19278__B1 _19207_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21469__B _21469_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14884__A2_N _22312_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12212_ _12190_/A _12210_/X _12211_/X VGND VGND VPWR VPWR _12212_/X sky130_fd_sc_hd__and3_4
X_15000_ _14879_/X _14982_/X _14880_/A VGND VGND VPWR VPWR _15001_/C sky130_fd_sc_hd__o21a_4
XFILLER_68_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13192_ _11711_/X _13173_/X _13191_/X _25001_/Q _13114_/X VGND VGND VPWR VPWR _13192_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__22821__A1 _21572_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25178_ _24847_/CLK _11822_/X HRESETn VGND VGND VPWR VPWR _25178_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12143_ _25106_/Q VGND VGND VPWR VPWR _12180_/B sky130_fd_sc_hd__inv_2
X_24129_ _24101_/CLK _16613_/X HRESETn VGND VGND VPWR VPWR _24129_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23741__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14269__A2_N _14268_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12074_ _12073_/Y _24576_/Q _12073_/Y _24576_/Q VGND VGND VPWR VPWR _12081_/B sky130_fd_sc_hd__a2bb2o_4
X_16951_ _16949_/Y _16950_/X _16951_/C VGND VGND VPWR VPWR _24062_/D sky130_fd_sc_hd__and3_4
XFILLER_123_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14899__A2_N _14897_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15902_ _24398_/Q VGND VGND VPWR VPWR _15902_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15483__A _15460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19670_ _23253_/Q VGND VGND VPWR VPWR _21910_/B sky130_fd_sc_hd__inv_2
X_16882_ _16881_/X VGND VGND VPWR VPWR _16882_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18621_ _18620_/Y VGND VGND VPWR VPWR _18621_/X sky130_fd_sc_hd__buf_2
X_15833_ _15826_/A VGND VGND VPWR VPWR _15847_/A sky130_fd_sc_hd__buf_2
XANTENNA__24947__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11516__A _16231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18552_ _18552_/A _18552_/B VGND VGND VPWR VPWR _18552_/X sky130_fd_sc_hd__or2_4
XFILLER_46_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19202__B1 _19201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15764_ _15748_/X _15763_/X _15600_/X _24452_/Q _15746_/X VGND VGND VPWR VPWR _15764_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12825__B1 _21840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12976_ _22308_/A _12976_/B VGND VGND VPWR VPWR _12976_/X sky130_fd_sc_hd__or2_4
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20829__A _21591_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17503_ _17503_/A _17503_/B VGND VGND VPWR VPWR _17515_/B sky130_fd_sc_hd__or2_4
XFILLER_45_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14715_ _14712_/X _14713_/Y _14997_/A _14714_/Y VGND VGND VPWR VPWR _14719_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20099__A2_N _20098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19753__B2 _19750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11927_ _21580_/A _11924_/X _25160_/Q _11924_/X VGND VGND VPWR VPWR _25161_/D sky130_fd_sc_hd__a2bb2o_4
X_18483_ _18483_/A VGND VGND VPWR VPWR _18483_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16567__A1 _15799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15695_ _15695_/A VGND VGND VPWR VPWR _15695_/X sky130_fd_sc_hd__buf_2
XFILLER_45_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17434_ _17323_/C _17408_/D VGND VGND VPWR VPWR _17434_/X sky130_fd_sc_hd__or2_4
X_14646_ _24727_/Q _14614_/B _24727_/Q _14614_/B VGND VGND VPWR VPWR _14646_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11858_ _11856_/Y _11852_/X _11857_/X _11852_/X VGND VGND VPWR VPWR _25170_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14837__A2_N _14835_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18050__A1_N _18049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17365_ _17362_/A _17358_/B _17364_/X VGND VGND VPWR VPWR _17365_/X sky130_fd_sc_hd__and3_4
X_11789_ _11772_/B _11786_/Y VGND VGND VPWR VPWR _11797_/A sky130_fd_sc_hd__and2_4
X_14577_ _17729_/A VGND VGND VPWR VPWR _14577_/X sky130_fd_sc_hd__buf_2
XFILLER_41_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19104_ _19103_/Y _19101_/X _19038_/X _19101_/X VGND VGND VPWR VPWR _23453_/D sky130_fd_sc_hd__a2bb2o_4
X_16316_ _24250_/Q VGND VGND VPWR VPWR _16316_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13528_ _13528_/A VGND VGND VPWR VPWR _13529_/B sky130_fd_sc_hd__inv_2
X_17296_ _17277_/X _17296_/B _17296_/C _17296_/D VGND VGND VPWR VPWR _17296_/X sky130_fd_sc_hd__or4_4
X_19035_ _19034_/Y VGND VGND VPWR VPWR _19035_/X sky130_fd_sc_hd__buf_2
X_16247_ _16247_/A VGND VGND VPWR VPWR _16247_/X sky130_fd_sc_hd__buf_2
XFILLER_9_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15658__A _15657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19269__B1 _19221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13459_ _16035_/A VGND VGND VPWR VPWR _13462_/A sky130_fd_sc_hd__inv_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23829__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21076__B1 _23618_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20037__A2_N _20036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16178_ _16196_/A VGND VGND VPWR VPWR _16178_/X sky130_fd_sc_hd__buf_2
XANTENNA__11564__B1 _11563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13178__A _13316_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15129_ _15129_/A _15123_/A _15117_/X VGND VGND VPWR VPWR _15130_/A sky130_fd_sc_hd__or3_4
XFILLER_47_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19937_ _21502_/B _19932_/X _19455_/A _19932_/X VGND VGND VPWR VPWR _23154_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15393__A _16376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19868_ _19868_/A VGND VGND VPWR VPWR _21780_/B sky130_fd_sc_hd__inv_2
XANTENNA__22040__A2 _22029_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16255__B1 _16254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24688__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18819_ _13194_/B VGND VGND VPWR VPWR _18819_/Y sky130_fd_sc_hd__inv_2
X_19799_ _19799_/A VGND VGND VPWR VPWR _19801_/A sky130_fd_sc_hd__buf_2
XFILLER_83_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22328__B1 _16658_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21830_ _22084_/A _20102_/Y VGND VGND VPWR VPWR _21830_/X sky130_fd_sc_hd__or2_4
XANTENNA__24617__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21842__B _22178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19744__B2 _19743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21761_ _21760_/X _19493_/Y VGND VGND VPWR VPWR _21761_/X sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_4_3_0_HCLK_A clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14737__A _14737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21551__B2 _21357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20712_ _20711_/X VGND VGND VPWR VPWR _23624_/D sky130_fd_sc_hd__inv_2
XANTENNA__24270__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23500_ _23560_/CLK _18976_/X VGND VGND VPWR VPWR _13123_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_23_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24480_ _24478_/CLK _24480_/D HRESETn VGND VGND VPWR VPWR _24480_/Q sky130_fd_sc_hd__dfrtp_4
X_21692_ _16042_/A _21691_/X _13622_/Y _22616_/A VGND VGND VPWR VPWR _21692_/X sky130_fd_sc_hd__o22a_4
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23431_ _23425_/CLK _19165_/X VGND VGND VPWR VPWR _17948_/B sky130_fd_sc_hd__dfxtp_4
X_20643_ _13524_/B VGND VGND VPWR VPWR _20643_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21303__B2 _21083_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23362_ _23350_/CLK _23362_/D VGND VGND VPWR VPWR _13210_/B sky130_fd_sc_hd__dfxtp_4
X_20574_ _20552_/X VGND VGND VPWR VPWR _20574_/X sky130_fd_sc_hd__buf_2
XANTENNA__17274__A1_N _25191_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18180__B1 _16054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22313_ _22226_/X _22312_/Y _16601_/Y _22228_/X VGND VGND VPWR VPWR _22313_/X sky130_fd_sc_hd__o22a_4
X_25101_ _23716_/CLK _12422_/X HRESETn VGND VGND VPWR VPWR _25101_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15568__A _11527_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23293_ _23293_/CLK _23293_/D VGND VGND VPWR VPWR _23293_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16730__B2 _22473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19285__A2_N _19284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12347__A2 _12346_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25032_ _24451_/CLK _12910_/X HRESETn VGND VGND VPWR VPWR _22900_/A sky130_fd_sc_hd__dfrtp_4
X_22244_ _22501_/A _22243_/X _21036_/X _24512_/Q _11530_/X VGND VGND VPWR VPWR _22245_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14741__B1 _14990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22803__A1 _24280_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13088__A _13011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12610__A2_N _24517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22175_ _22175_/A _22175_/B _22172_/X _22174_/X VGND VGND VPWR VPWR _22182_/A sky130_fd_sc_hd__or4_4
XANTENNA__16494__B1 _15479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20290__A1 _14234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21126_ _13334_/X _21066_/B _21126_/C VGND VGND VPWR VPWR _21127_/D sky130_fd_sc_hd__and3_4
XFILLER_120_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21057_ _21432_/C VGND VGND VPWR VPWR _22835_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_115_0_HCLK clkbuf_7_57_0_HCLK/X VGND VGND VPWR VPWR _24879_/CLK sky130_fd_sc_hd__clkbuf_1
X_20008_ _20007_/Y _20003_/X _15416_/X _19990_/Y VGND VGND VPWR VPWR _23127_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_178_0_HCLK clkbuf_7_89_0_HCLK/X VGND VGND VPWR VPWR _24521_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__17994__B1 _23917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22848__B _13618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12830_ _12829_/Y VGND VGND VPWR VPWR _12964_/A sky130_fd_sc_hd__buf_2
XANTENNA__24358__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24816_ _23774_/CLK _14222_/X HRESETn VGND VGND VPWR VPWR _20336_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_76_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12761_ _12761_/A VGND VGND VPWR VPWR _25041_/D sky130_fd_sc_hd__inv_2
XPHY_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24747_ _24748_/CLK _14520_/X HRESETn VGND VGND VPWR VPWR _21752_/A sky130_fd_sc_hd__dfrtp_4
X_21959_ _21955_/X _21958_/X _14524_/D VGND VGND VPWR VPWR _21959_/Y sky130_fd_sc_hd__o21ai_4
XPHY_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _24749_/Q VGND VGND VPWR VPWR _14500_/Y sky130_fd_sc_hd__inv_2
X_11712_ _18638_/A _18638_/B _11711_/X VGND VGND VPWR VPWR _11712_/X sky130_fd_sc_hd__o21a_4
XFILLER_70_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12677_/X VGND VGND VPWR VPWR _12692_/Y sky130_fd_sc_hd__inv_2
X_15480_ _15368_/X _15461_/X _15479_/X _24570_/Q _15466_/X VGND VGND VPWR VPWR _24570_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24678_ _24681_/CLK _15135_/Y HRESETn VGND VGND VPWR VPWR _24678_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22864__A _22351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11643_/A VGND VGND VPWR VPWR _11643_/X sky130_fd_sc_hd__buf_2
X_14431_ _14431_/A VGND VGND VPWR VPWR _14435_/B sky130_fd_sc_hd__inv_2
XFILLER_30_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23629_ _23648_/CLK _20276_/Y HRESETn VGND VGND VPWR VPWR _23629_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12167__A _24500_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17150_ _17144_/A _17153_/B VGND VGND VPWR VPWR _17150_/Y sky130_fd_sc_hd__nand2_4
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11574_ _11572_/Y _11569_/X _11573_/X _11569_/X VGND VGND VPWR VPWR _25207_/D sky130_fd_sc_hd__a2bb2o_4
X_14362_ _14362_/A VGND VGND VPWR VPWR _14362_/Y sky130_fd_sc_hd__inv_2
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23993__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16101_ _16098_/Y _16099_/X _16100_/X _16099_/X VGND VGND VPWR VPWR _16101_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13313_ _13137_/A _13313_/B VGND VGND VPWR VPWR _13314_/C sky130_fd_sc_hd__or2_4
XFILLER_128_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14293_ _14288_/A VGND VGND VPWR VPWR _14293_/X sky130_fd_sc_hd__buf_2
X_17081_ _17026_/A _17079_/A VGND VGND VPWR VPWR _17081_/X sky130_fd_sc_hd__or2_4
XANTENNA__23922__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25146__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13244_ _13244_/A _23473_/Q VGND VGND VPWR VPWR _13244_/X sky130_fd_sc_hd__or2_4
X_16032_ _16032_/A VGND VGND VPWR VPWR _16032_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11546__B1 _11545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13175_ _13137_/A _13175_/B VGND VGND VPWR VPWR _13175_/X sky130_fd_sc_hd__or2_4
XFILLER_123_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12126_ _12299_/A _12124_/Y _12122_/A _12125_/Y VGND VGND VPWR VPWR _12131_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11561__A3 HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17983_ _17974_/X VGND VGND VPWR VPWR _17983_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_11_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_97_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19722_ _19720_/Y _19718_/X _19721_/X _19718_/X VGND VGND VPWR VPWR _19722_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_74_0_HCLK clkbuf_7_74_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_74_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12057_ _12011_/Y _12056_/Y SCLK_S3 _12055_/X VGND VGND VPWR VPWR _12057_/X sky130_fd_sc_hd__o22a_4
X_16934_ _16936_/A _16927_/X _16934_/C VGND VGND VPWR VPWR _16934_/X sky130_fd_sc_hd__and3_4
XFILLER_96_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19653_ _21832_/B _19647_/X _19603_/X _19652_/X VGND VGND VPWR VPWR _19653_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24781__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16865_ _24086_/Q _16864_/Y VGND VGND VPWR VPWR _16867_/B sky130_fd_sc_hd__or2_4
XFILLER_37_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17985__B1 _15501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18604_ _18561_/Y _18482_/A _18582_/X _18603_/X VGND VGND VPWR VPWR _18604_/X sky130_fd_sc_hd__o22a_4
XFILLER_92_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15816_ _15712_/X _15815_/Y _15713_/X _15815_/Y VGND VGND VPWR VPWR _15816_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14799__B1 _15045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24099__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24710__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19584_ _21674_/B _19581_/X _19452_/X _19581_/X VGND VGND VPWR VPWR _23283_/D sky130_fd_sc_hd__a2bb2o_4
X_16796_ _16792_/X _16793_/X _16796_/C _16795_/X VGND VGND VPWR VPWR _16796_/X sky130_fd_sc_hd__or4_4
XFILLER_65_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18535_ _18535_/A _18535_/B VGND VGND VPWR VPWR _18536_/B sky130_fd_sc_hd__or2_4
XFILLER_0_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24028__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15747_ _15693_/X _15740_/X _15743_/X _24460_/Q _15746_/X VGND VGND VPWR VPWR _24460_/D
+ sky130_fd_sc_hd__a32o_4
X_12959_ _12952_/A _12959_/B _12958_/X VGND VGND VPWR VPWR _12959_/X sky130_fd_sc_hd__and3_4
XANTENNA__13461__A _11507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21533__B2 _21400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18466_ _18482_/A _18466_/B _18465_/X VGND VGND VPWR VPWR _18467_/A sky130_fd_sc_hd__or3_4
X_15678_ _12319_/Y _15677_/X _15350_/X _15677_/X VGND VGND VPWR VPWR _15678_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17417_ _17319_/Y _17419_/B _17416_/Y VGND VGND VPWR VPWR _17417_/X sky130_fd_sc_hd__o21a_4
XFILLER_18_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14629_ _14628_/X VGND VGND VPWR VPWR _14630_/B sky130_fd_sc_hd__inv_2
X_18397_ _23833_/Q VGND VGND VPWR VPWR _18488_/A sky130_fd_sc_hd__inv_2
XANTENNA__16960__B2 _24058_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17348_ _17303_/Y _17348_/B _17288_/Y _17348_/D VGND VGND VPWR VPWR _17349_/B sky130_fd_sc_hd__or4_4
XFILLER_119_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17279_ _11554_/Y _24001_/Q _11554_/Y _24001_/Q VGND VGND VPWR VPWR _17279_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12805__A _22133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19018_ _19012_/Y VGND VGND VPWR VPWR _19018_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20290_ _14234_/Y _20273_/X _20287_/X _20289_/X VGND VGND VPWR VPWR _20291_/A sky130_fd_sc_hd__a211o_4
XFILLER_127_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22797__B1 _22178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21903__A2_N _22153_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22013__A2 _20749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19414__B1 _19392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22204__A1_N _12345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23980_ _25194_/CLK _17440_/X HRESETn VGND VGND VPWR VPWR _17264_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_29_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22931_ _22931_/A _22928_/X _22930_/X VGND VGND VPWR VPWR _22931_/X sky130_fd_sc_hd__and3_4
XANTENNA__16779__A1 _24397_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15851__A _24417_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24451__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21572__B _21572_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22862_ _22334_/A _22862_/B _22862_/C VGND VGND VPWR VPWR _22874_/B sky130_fd_sc_hd__and3_4
X_24601_ _24604_/CLK _15362_/X HRESETn VGND VGND VPWR VPWR _15361_/A sky130_fd_sc_hd__dfrtp_4
X_21813_ _20962_/A _21811_/X _21812_/X VGND VGND VPWR VPWR _21813_/X sky130_fd_sc_hd__and3_4
XANTENNA__17991__A3 _16451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22793_ _16325_/Y _20757_/A _16063_/Y _22548_/A VGND VGND VPWR VPWR _22793_/X sky130_fd_sc_hd__o22a_4
X_21744_ _21079_/X _21738_/Y _21308_/X _21743_/X VGND VGND VPWR VPWR _21744_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24532_ _24478_/CLK _15587_/X HRESETn VGND VGND VPWR VPWR _24532_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21675_ _21675_/A _21675_/B _21674_/X VGND VGND VPWR VPWR _21675_/X sky130_fd_sc_hd__and3_4
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24463_ _24944_/CLK _15737_/X HRESETn VGND VGND VPWR VPWR _20738_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_12_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20626_ _20635_/C _13537_/C VGND VGND VPWR VPWR _20627_/A sky130_fd_sc_hd__or2_4
XFILLER_32_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23414_ _25194_/CLK _19214_/X VGND VGND VPWR VPWR _22046_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24394_ _24071_/CLK _24394_/D HRESETn VGND VGND VPWR VPWR _20737_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_137_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23345_ _23336_/CLK _23345_/D VGND VGND VPWR VPWR _13249_/B sky130_fd_sc_hd__dfxtp_4
X_20557_ _16555_/Y _20553_/X _13526_/B _20556_/X VGND VGND VPWR VPWR _20558_/A sky130_fd_sc_hd__o22a_4
XANTENNA__16703__A1 _22783_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23276_ _23258_/CLK _23276_/D VGND VGND VPWR VPWR _23276_/Q sky130_fd_sc_hd__dfxtp_4
X_20488_ _20465_/A VGND VGND VPWR VPWR _20488_/X sky130_fd_sc_hd__buf_2
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22227_ _14923_/Y _22227_/B VGND VGND VPWR VPWR _22227_/X sky130_fd_sc_hd__and2_4
XFILLER_4_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25015_ _25034_/CLK _25015_/D HRESETn VGND VGND VPWR VPWR _22258_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_106_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23665__D _23665_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14854__A1_N _14712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22158_ _21050_/Y VGND VGND VPWR VPWR _22163_/A sky130_fd_sc_hd__buf_2
XFILLER_43_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21109_ _15403_/Y _21109_/B VGND VGND VPWR VPWR _21109_/X sky130_fd_sc_hd__and2_4
XANTENNA__19405__B1 _19381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24539__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14980_ _14697_/Y _14980_/B VGND VGND VPWR VPWR _14981_/C sky130_fd_sc_hd__or2_4
X_22089_ _22089_/A _22089_/B _22088_/X VGND VGND VPWR VPWR _22089_/X sky130_fd_sc_hd__and3_4
XFILLER_102_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22859__A _22859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13931_ _13930_/X VGND VGND VPWR VPWR _13931_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15761__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24192__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16650_ _16643_/A VGND VGND VPWR VPWR _16650_/X sky130_fd_sc_hd__buf_2
X_13862_ _13862_/A VGND VGND VPWR VPWR _13862_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15442__A1 RsRx_S0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15601_ _15574_/X _15599_/X _15600_/X _24525_/Q _15585_/X VGND VGND VPWR VPWR _15601_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24121__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12813_ _12813_/A VGND VGND VPWR VPWR _12813_/Y sky130_fd_sc_hd__inv_2
X_16581_ _16581_/A VGND VGND VPWR VPWR _16581_/X sky130_fd_sc_hd__buf_2
XFILLER_62_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13793_ _13794_/A _13793_/B VGND VGND VPWR VPWR _13793_/X sky130_fd_sc_hd__and2_4
XFILLER_103_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18320_ _18303_/X _18320_/B _18319_/X VGND VGND VPWR VPWR _18320_/X sky130_fd_sc_hd__and3_4
X_15532_ _15430_/X _15319_/Y _15432_/X _13519_/A _15531_/X VGND VGND VPWR VPWR _15532_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_103_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12744_ _12649_/C _12747_/B _12666_/X VGND VGND VPWR VPWR _12744_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__17195__A1 _23766_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22594__A _21051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18251_ _18242_/A _18250_/X _18228_/X VGND VGND VPWR VPWR _18251_/Y sky130_fd_sc_hd__a21oi_4
X_15463_ _15463_/A VGND VGND VPWR VPWR _15463_/X sky130_fd_sc_hd__buf_2
X_12675_ _12669_/A _12663_/X _12674_/X _12671_/B VGND VGND VPWR VPWR _12676_/A sky130_fd_sc_hd__a211o_4
XFILLER_31_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17202_ _16373_/A VGND VGND VPWR VPWR _17202_/X sky130_fd_sc_hd__buf_2
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ _14414_/A _14378_/A VGND VGND VPWR VPWR _14414_/X sky130_fd_sc_hd__or2_4
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _13632_/A VGND VGND VPWR VPWR _11626_/X sky130_fd_sc_hd__buf_2
X_18182_ _16058_/Y _23871_/Q _24344_/Q _18207_/B VGND VGND VPWR VPWR _18182_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22744__D _22743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15394_ _21728_/A _15387_/X _15393_/X _15387_/X VGND VGND VPWR VPWR _24589_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ _17133_/A _17133_/B VGND VGND VPWR VPWR _17154_/A sky130_fd_sc_hd__or2_4
XFILLER_128_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ _14335_/X _14344_/X _24785_/Q _14320_/Y VGND VGND VPWR VPWR _14345_/X sky130_fd_sc_hd__o22a_4
X_11557_ _25212_/Q VGND VGND VPWR VPWR _11557_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22491__A2 _22173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17064_ _17052_/A _17064_/B _17064_/C VGND VGND VPWR VPWR _17064_/X sky130_fd_sc_hd__and3_4
XANTENNA__21938__A _21339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14276_ _14275_/Y _14273_/X _14209_/X _14273_/X VGND VGND VPWR VPWR _14276_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20842__A _16043_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16015_ _16221_/C _16012_/X _24359_/Q _16014_/X VGND VGND VPWR VPWR _16015_/X sky130_fd_sc_hd__o22a_4
X_13227_ _13120_/X _13227_/B VGND VGND VPWR VPWR _13227_/X sky130_fd_sc_hd__or2_4
XFILLER_98_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16458__B1 _16369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24962__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13158_ _13122_/A _13156_/X _13157_/X VGND VGND VPWR VPWR _13158_/X sky130_fd_sc_hd__and3_4
XFILLER_124_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12109_ _25131_/Q _24574_/Q _12170_/A _12108_/Y VGND VGND VPWR VPWR _12119_/A sky130_fd_sc_hd__o22a_4
X_13089_ _11733_/A VGND VGND VPWR VPWR _13247_/A sky130_fd_sc_hd__buf_2
X_17966_ _17934_/A _17966_/B VGND VGND VPWR VPWR _17968_/B sky130_fd_sc_hd__or2_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16917_ _16936_/A _16917_/B _16917_/C VGND VGND VPWR VPWR _24072_/D sky130_fd_sc_hd__and3_4
X_19705_ _23239_/Q VGND VGND VPWR VPWR _20972_/B sky130_fd_sc_hd__inv_2
XANTENNA__24209__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17897_ _17929_/A _17895_/X _17897_/C VGND VGND VPWR VPWR _17898_/C sky130_fd_sc_hd__and3_4
XFILLER_38_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22488__B _22488_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16848_ _16940_/A VGND VGND VPWR VPWR _16858_/A sky130_fd_sc_hd__inv_2
X_19636_ _19636_/A VGND VGND VPWR VPWR _19636_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_161_0_HCLK clkbuf_7_80_0_HCLK/X VGND VGND VPWR VPWR _23493_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_4_0_HCLK clkbuf_7_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_4_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16630__B1 HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19567_ _19554_/Y VGND VGND VPWR VPWR _19567_/X sky130_fd_sc_hd__buf_2
XFILLER_65_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_18_0_HCLK clkbuf_7_9_0_HCLK/X VGND VGND VPWR VPWR _23898_/CLK sky130_fd_sc_hd__clkbuf_1
X_16779_ _24397_/Q _24061_/Q _15904_/Y _16778_/Y VGND VGND VPWR VPWR _16782_/C sky130_fd_sc_hd__o22a_4
XFILLER_94_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14287__A _16559_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18982__A _18982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18518_ _18518_/A _18518_/B VGND VGND VPWR VPWR _18519_/C sky130_fd_sc_hd__or2_4
XFILLER_59_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19498_ _23314_/Q VGND VGND VPWR VPWR _19498_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18449_ _18475_/A VGND VGND VPWR VPWR _18449_/X sky130_fd_sc_hd__buf_2
XANTENNA__17598__A _17595_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23844__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12012__A1_N _12011_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25068__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21460_ _21935_/A _21460_/B VGND VGND VPWR VPWR _21461_/C sky130_fd_sc_hd__or2_4
XANTENNA__14734__B _14727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20411_ _20227_/A _20232_/C _15250_/X VGND VGND VPWR VPWR _23687_/D sky130_fd_sc_hd__o21a_4
X_21391_ _21387_/A _21391_/B _21390_/X VGND VGND VPWR VPWR _21391_/X sky130_fd_sc_hd__and3_4
XFILLER_88_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23130_ _23128_/CLK _23130_/D VGND VGND VPWR VPWR _20000_/A sky130_fd_sc_hd__dfxtp_4
X_20342_ _13794_/A _15250_/X _13790_/X VGND VGND VPWR VPWR _20342_/X sky130_fd_sc_hd__and3_4
XANTENNA__20752__A _20751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23061_ _20739_/X VGND VGND VPWR VPWR IRQ[9] sky130_fd_sc_hd__buf_2
X_20273_ _20296_/A VGND VGND VPWR VPWR _20273_/X sky130_fd_sc_hd__buf_2
XANTENNA__21567__B _22445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22012_ _16537_/Y _20866_/A VGND VGND VPWR VPWR _22012_/X sky130_fd_sc_hd__and2_4
XFILLER_89_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16449__B1 _16279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21583__A _13324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23963_ _23949_/CLK _17555_/X HRESETn VGND VGND VPWR VPWR _16692_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_99_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21745__A1 _21564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22398__B _22395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22914_ _23026_/B _22913_/X _22459_/X _24530_/Q _22460_/X VGND VGND VPWR VPWR _22914_/X
+ sky130_fd_sc_hd__a32o_4
X_23894_ _24748_/CLK _18078_/X HRESETn VGND VGND VPWR VPWR _23894_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19988__A _23134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22845_ _23026_/B _22844_/X _22459_/X _24528_/Q _22460_/X VGND VGND VPWR VPWR _22845_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14197__A _14197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11614__A _11614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22776_ _16413_/Y _22551_/X _14729_/Y _22547_/X VGND VGND VPWR VPWR _22777_/B sky130_fd_sc_hd__o22a_4
XANTENNA__20927__A _20926_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24515_ _24483_/CLK _24515_/D HRESETn VGND VGND VPWR VPWR _24515_/Q sky130_fd_sc_hd__dfrtp_4
X_21727_ _20575_/Y _21280_/X _20438_/Y _21562_/A VGND VGND VPWR VPWR _21727_/X sky130_fd_sc_hd__o22a_4
XFILLER_40_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12460_ _12460_/A _12448_/B _12459_/X VGND VGND VPWR VPWR _12460_/X sky130_fd_sc_hd__and3_4
X_21658_ _21009_/A VGND VGND VPWR VPWR _21677_/A sky130_fd_sc_hd__buf_2
XFILLER_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24446_ _24445_/CLK _24446_/D HRESETn VGND VGND VPWR VPWR _24446_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12391_ _12391_/A VGND VGND VPWR VPWR _12391_/Y sky130_fd_sc_hd__inv_2
X_20609_ _20611_/A VGND VGND VPWR VPWR _20609_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21589_ _12001_/Y _22840_/A _21587_/X _21881_/A VGND VGND VPWR VPWR _21600_/B sky130_fd_sc_hd__a211o_4
XANTENNA__19874__B1 _19828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24377_ _24385_/CLK _15958_/X HRESETn VGND VGND VPWR VPWR _15957_/A sky130_fd_sc_hd__dfrtp_4
X_14130_ _24847_/Q _14122_/X _24846_/Q _14127_/X VGND VGND VPWR VPWR _14130_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21758__A _15572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23328_ _23135_/CLK _23328_/D VGND VGND VPWR VPWR _19461_/A sky130_fd_sc_hd__dfxtp_4
X_14061_ _14059_/Y _14060_/X _13638_/X _14060_/X VGND VGND VPWR VPWR _24866_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15360__B1 _11570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15756__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23259_ _23258_/CLK _23259_/D VGND VGND VPWR VPWR _19654_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__20236__A1 _24822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13012_ _11743_/A VGND VGND VPWR VPWR _13045_/A sky130_fd_sc_hd__buf_2
XANTENNA__21433__B1 _21107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_6_0_HCLK_A clkbuf_5_6_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17820_ _17721_/A VGND VGND VPWR VPWR _17821_/A sky130_fd_sc_hd__buf_2
XANTENNA__13276__A _13182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24373__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22589__A _22588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17751_ _17676_/X _17751_/B _17750_/X VGND VGND VPWR VPWR _17752_/C sky130_fd_sc_hd__and3_4
XFILLER_88_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24302__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14963_ _14954_/X _14957_/X _14959_/X _14962_/X VGND VGND VPWR VPWR _14973_/C sky130_fd_sc_hd__or4_4
XANTENNA__13674__B1 _13398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21736__B2 _21425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21997__A1_N _20747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25186__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16702_ _22782_/A VGND VGND VPWR VPWR _16702_/Y sky130_fd_sc_hd__inv_2
X_13914_ _24899_/Q _13908_/X _13905_/X _13810_/X _13911_/X VGND VGND VPWR VPWR _13914_/X
+ sky130_fd_sc_hd__a32o_4
X_17682_ _17698_/A _17682_/B VGND VGND VPWR VPWR _17682_/X sky130_fd_sc_hd__or2_4
XFILLER_74_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14894_ _14894_/A VGND VGND VPWR VPWR _14895_/A sky130_fd_sc_hd__inv_2
XFILLER_63_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19421_ HWDATA[6] VGND VGND VPWR VPWR _19421_/X sky130_fd_sc_hd__buf_2
XFILLER_90_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16612__B1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16633_ _14714_/Y _16629_/X HWDATA[27] _16632_/X VGND VGND VPWR VPWR _24120_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_234_0_HCLK clkbuf_8_235_0_HCLK/A VGND VGND VPWR VPWR _25097_/CLK sky130_fd_sc_hd__clkbuf_1
X_13845_ _13845_/A _13806_/X _13811_/C _13810_/X VGND VGND VPWR VPWR _13845_/X sky130_fd_sc_hd__or4_4
X_19352_ _23365_/Q VGND VGND VPWR VPWR _19352_/Y sky130_fd_sc_hd__inv_2
X_16564_ _23008_/B VGND VGND VPWR VPWR _22228_/A sky130_fd_sc_hd__buf_2
X_13776_ _13764_/X _13776_/B _13776_/C _13775_/Y VGND VGND VPWR VPWR _13777_/D sky130_fd_sc_hd__and4_4
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20837__A _20800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18303_ _18318_/A _18302_/X VGND VGND VPWR VPWR _18303_/X sky130_fd_sc_hd__or2_4
XFILLER_71_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15515_ _12098_/Y _15509_/X _15513_/X _15514_/X VGND VGND VPWR VPWR _15515_/X sky130_fd_sc_hd__a2bb2o_4
X_12727_ _12727_/A _12653_/C VGND VGND VPWR VPWR _12728_/B sky130_fd_sc_hd__or2_4
X_19283_ _19283_/A VGND VGND VPWR VPWR _19283_/Y sky130_fd_sc_hd__inv_2
X_16495_ _16495_/A VGND VGND VPWR VPWR _16495_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14835__A _24129_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25161__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18234_ _18234_/A _18234_/B VGND VGND VPWR VPWR _18236_/B sky130_fd_sc_hd__or2_4
X_15446_ _15438_/A _15437_/X _15449_/B _14434_/A _15445_/Y VGND VGND VPWR VPWR _24580_/D
+ sky130_fd_sc_hd__a32o_4
X_12658_ _12657_/X VGND VGND VPWR VPWR _12658_/Y sky130_fd_sc_hd__inv_2
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11609_ _25197_/Q VGND VGND VPWR VPWR _11609_/Y sky130_fd_sc_hd__inv_2
X_18165_ _23862_/Q VGND VGND VPWR VPWR _18278_/A sky130_fd_sc_hd__inv_2
XFILLER_129_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15377_ _22323_/A _15374_/X _11598_/X _15374_/X VGND VGND VPWR VPWR _24595_/D sky130_fd_sc_hd__a2bb2o_4
X_12589_ _25055_/Q _12588_/A _12587_/Y _12588_/Y VGND VGND VPWR VPWR _12590_/D sky130_fd_sc_hd__o22a_4
XFILLER_50_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17116_ _17116_/A _17116_/B VGND VGND VPWR VPWR _17116_/X sky130_fd_sc_hd__or2_4
XFILLER_8_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16679__B1 _16678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14328_ _24780_/Q _14325_/X _14326_/Y _14327_/X VGND VGND VPWR VPWR _14329_/B sky130_fd_sc_hd__o22a_4
X_18096_ _18095_/X VGND VGND VPWR VPWR _18096_/Y sky130_fd_sc_hd__inv_2
X_17047_ _17070_/A _17046_/X VGND VGND VPWR VPWR _17054_/A sky130_fd_sc_hd__or2_4
XANTENNA__15351__B1 _15350_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14259_ _14259_/A VGND VGND VPWR VPWR _14259_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21975__B2 _21187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13186__A _11741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18998_ _23491_/Q VGND VGND VPWR VPWR _21655_/B sky130_fd_sc_hd__inv_2
XFILLER_135_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22519__A3 _21981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24043__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_44_0_HCLK clkbuf_6_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_44_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17949_ _17853_/A _17949_/B VGND VGND VPWR VPWR _17950_/C sky130_fd_sc_hd__or2_4
XFILLER_26_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21727__B2 _21562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20960_ _20965_/A VGND VGND VPWR VPWR _20961_/A sky130_fd_sc_hd__buf_2
XFILLER_66_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16603__B1 _15507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19619_ _19619_/A VGND VGND VPWR VPWR _20966_/B sky130_fd_sc_hd__inv_2
X_20891_ _20891_/A _13326_/A VGND VGND VPWR VPWR _20891_/X sky130_fd_sc_hd__or2_4
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22630_ _22116_/X _22628_/X _22629_/X _24564_/Q _22118_/X VGND VGND VPWR VPWR _22631_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_59_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22152__A1 _22879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20747__A _15821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11979__B1 _11636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22152__B2 _22151_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22561_ _24412_/Q _22557_/X _22558_/X _22560_/X VGND VGND VPWR VPWR _22562_/C sky130_fd_sc_hd__a211o_4
XANTENNA__16252__A1_N _14913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21512_ _14471_/A _21512_/B _21511_/X VGND VGND VPWR VPWR _21512_/X sky130_fd_sc_hd__or3_4
X_24300_ _24319_/CLK _24300_/D HRESETn VGND VGND VPWR VPWR _24300_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22492_ _16436_/Y _21882_/X _16649_/Y _22017_/X VGND VGND VPWR VPWR _22492_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21443_ _21443_/A _21097_/B VGND VGND VPWR VPWR _21443_/X sky130_fd_sc_hd__and2_4
X_24231_ _23840_/CLK _16365_/X HRESETn VGND VGND VPWR VPWR _16363_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_21_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16267__A1_N _14933_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24162_ _24162_/CLK _16547_/X HRESETn VGND VGND VPWR VPWR _16544_/A sky130_fd_sc_hd__dfrtp_4
X_21374_ _21374_/A _21374_/B VGND VGND VPWR VPWR _21374_/X sky130_fd_sc_hd__or2_4
XFILLER_108_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24884__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20325_ _13921_/A _20322_/X _20324_/X VGND VGND VPWR VPWR _23640_/D sky130_fd_sc_hd__and3_4
XFILLER_107_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15576__A _15575_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23113_ _23293_/CLK _20046_/X VGND VGND VPWR VPWR _23113_/Q sky130_fd_sc_hd__dfxtp_4
X_24093_ _24094_/CLK _24093_/D HRESETn VGND VGND VPWR VPWR _24093_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14480__A _14480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21415__B1 _24505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_126_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_253_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_23044_ VGND VGND VPWR VPWR _23044_/HI IRQ[12] sky130_fd_sc_hd__conb_1
X_20256_ _23770_/Q _20225_/B _20224_/B _20255_/Y VGND VGND VPWR VPWR _20257_/D sky130_fd_sc_hd__a211o_4
XANTENNA__20769__A2 _20765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13096__A _11741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11609__A _25197_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20187_ _20173_/A _20185_/Y VGND VGND VPWR VPWR _20187_/X sky130_fd_sc_hd__or2_4
XFILLER_44_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13656__B1 _11598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22202__A _22202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24995_ _25159_/CLK _13331_/X HRESETn VGND VGND VPWR VPWR _23041_/A sky130_fd_sc_hd__dfrtp_4
X_11960_ _11960_/A VGND VGND VPWR VPWR _13333_/A sky130_fd_sc_hd__buf_2
X_23946_ _23972_/CLK _23946_/D HRESETn VGND VGND VPWR VPWR _23946_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18595__B1 _16351_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13543__B _13543_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11891_ _11891_/A VGND VGND VPWR VPWR _11891_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23766__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23877_ _24088_/CLK _23877_/D HRESETn VGND VGND VPWR VPWR _20736_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__22856__B _22853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13630_ _16043_/A _23763_/Q _13630_/C _22314_/B VGND VGND VPWR VPWR _13630_/X sky130_fd_sc_hd__and4_4
XFILLER_32_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22828_ _17482_/A _22654_/X _22608_/X VGND VGND VPWR VPWR _22830_/C sky130_fd_sc_hd__a21o_4
XANTENNA__22143__A1 _21564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21734__A2_N _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22143__B2 _22142_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_64_0_HCLK clkbuf_8_65_0_HCLK/A VGND VGND VPWR VPWR _24851_/CLK sky130_fd_sc_hd__clkbuf_1
X_13561_ _11679_/Y _13561_/B VGND VGND VPWR VPWR _13562_/B sky130_fd_sc_hd__or2_4
XFILLER_73_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22694__A2 _21553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22759_ _22681_/A _22759_/B VGND VGND VPWR VPWR _22759_/X sky130_fd_sc_hd__and2_4
X_15300_ _23762_/D VGND VGND VPWR VPWR _15300_/Y sky130_fd_sc_hd__inv_2
X_12512_ _12406_/Y _12511_/X _12444_/A _12507_/B VGND VGND VPWR VPWR _12512_/X sky130_fd_sc_hd__a211o_4
XFILLER_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16280_ _14897_/Y _16278_/X _16279_/X _16278_/X VGND VGND VPWR VPWR _16280_/X sky130_fd_sc_hd__a2bb2o_4
X_13492_ _13492_/A VGND VGND VPWR VPWR _13492_/X sky130_fd_sc_hd__buf_2
XFILLER_100_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15231_ _15222_/X _15231_/B _15226_/C VGND VGND VPWR VPWR _24651_/D sky130_fd_sc_hd__and3_4
X_12443_ _12415_/X _12424_/B _12416_/A VGND VGND VPWR VPWR _12443_/X sky130_fd_sc_hd__o21a_4
X_24429_ _24432_/CLK _24429_/D HRESETn VGND VGND VPWR VPWR _20834_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22446__A2 _22227_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12395__B1 _12389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15162_ _15162_/A VGND VGND VPWR VPWR _15163_/B sky130_fd_sc_hd__inv_2
XFILLER_125_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21488__A _17636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12374_ _12411_/A VGND VGND VPWR VPWR _12489_/A sky130_fd_sc_hd__buf_2
XANTENNA__17685__B _17685_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14113_ _24852_/Q _14112_/Y _14106_/B VGND VGND VPWR VPWR _24852_/D sky130_fd_sc_hd__o21a_4
XFILLER_4_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24554__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15093_ _14867_/A _15093_/B _15093_/C VGND VGND VPWR VPWR _15093_/X sky130_fd_sc_hd__and3_4
X_19970_ _19982_/A VGND VGND VPWR VPWR _19970_/X sky130_fd_sc_hd__buf_2
XANTENNA__12903__A _12921_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21406__B1 _21793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14044_ _14043_/Y _14027_/X _13635_/X _14027_/X VGND VGND VPWR VPWR _24872_/D sky130_fd_sc_hd__a2bb2o_4
X_18921_ _18920_/X VGND VGND VPWR VPWR _18935_/A sky130_fd_sc_hd__inv_2
XFILLER_4_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18852_ _18968_/A _18072_/X _18069_/X VGND VGND VPWR VPWR _18852_/X sky130_fd_sc_hd__or3_4
XFILLER_95_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21935__B _21935_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15636__A1 _15619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15636__B2 _15585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17803_ _17689_/X _17803_/B _17802_/X VGND VGND VPWR VPWR _17803_/X sky130_fd_sc_hd__and3_4
XFILLER_94_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18783_ _18920_/A _19123_/B _14587_/X _19123_/D VGND VGND VPWR VPWR _18784_/A sky130_fd_sc_hd__or4_4
X_15995_ _24363_/Q VGND VGND VPWR VPWR _15995_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22112__A _20968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17734_ _17781_/A _23421_/Q VGND VGND VPWR VPWR _17737_/B sky130_fd_sc_hd__or2_4
XFILLER_94_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14946_ _24673_/Q VGND VGND VPWR VPWR _14946_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21951__A _21394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17665_ _17662_/B _17655_/X VGND VGND VPWR VPWR _17665_/X sky130_fd_sc_hd__or2_4
XFILLER_78_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14877_ _14762_/Y _14757_/Y _14875_/X _14877_/D VGND VGND VPWR VPWR _14877_/X sky130_fd_sc_hd__or4_4
XFILLER_78_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20932__A2 _11940_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16616_ _24126_/Q VGND VGND VPWR VPWR _16616_/Y sky130_fd_sc_hd__inv_2
X_19404_ _19404_/A VGND VGND VPWR VPWR _19404_/Y sky130_fd_sc_hd__inv_2
X_13828_ _13828_/A _13816_/A _13828_/C _13828_/D VGND VGND VPWR VPWR _13831_/C sky130_fd_sc_hd__or4_4
XANTENNA__16600__A3 _16096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19421__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17596_ _17490_/A _17595_/X _17528_/X _17591_/B VGND VGND VPWR VPWR _17597_/A sky130_fd_sc_hd__a211o_4
XFILLER_1_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16547_ _16544_/Y _16542_/X _16546_/X _16542_/X VGND VGND VPWR VPWR _16547_/X sky130_fd_sc_hd__a2bb2o_4
X_19335_ _19333_/Y _19328_/X _19311_/X _19334_/X VGND VGND VPWR VPWR _19335_/X sky130_fd_sc_hd__a2bb2o_4
X_13759_ _13753_/A VGND VGND VPWR VPWR _13776_/B sky130_fd_sc_hd__inv_2
XFILLER_56_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19266_ _19260_/X VGND VGND VPWR VPWR _19266_/X sky130_fd_sc_hd__buf_2
XANTENNA__21893__B1 _23622_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12395__A2_N _24473_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16478_ _16475_/X VGND VGND VPWR VPWR _16479_/A sky130_fd_sc_hd__inv_2
XANTENNA__22782__A _22782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18217_ _18210_/X _18213_/X _18217_/C VGND VGND VPWR VPWR _18218_/C sky130_fd_sc_hd__or3_4
X_15429_ _15428_/X VGND VGND VPWR VPWR _15430_/A sky130_fd_sc_hd__buf_2
X_19197_ _19195_/Y _19191_/X _19152_/X _19196_/X VGND VGND VPWR VPWR _19197_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22437__A2 _22435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12085__A _24555_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18148_ _23853_/Q VGND VGND VPWR VPWR _18210_/B sky130_fd_sc_hd__inv_2
XANTENNA__17595__B _16700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15396__A _15401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24295__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18079_ _21188_/A _18065_/B _11765_/A VGND VGND VPWR VPWR _18080_/A sky130_fd_sc_hd__o21a_4
XFILLER_102_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20110_ _20110_/A VGND VGND VPWR VPWR _20110_/X sky130_fd_sc_hd__buf_2
XANTENNA__24224__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21090_ _21082_/X _21090_/B _21087_/X _21090_/D VGND VGND VPWR VPWR _21090_/X sky130_fd_sc_hd__or4_4
XFILLER_131_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20041_ _20035_/Y VGND VGND VPWR VPWR _20041_/X sky130_fd_sc_hd__buf_2
XFILLER_59_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23763__D _20197_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13644__A _13644_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23800_ _23796_/CLK _12045_/C HRESETn VGND VGND VPWR VPWR _12040_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_22_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19561__A2_N _19555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24780_ _23618_/CLK _14329_/X HRESETn VGND VGND VPWR VPWR _24780_/Q sky130_fd_sc_hd__dfrtp_4
X_21992_ _22249_/A VGND VGND VPWR VPWR _22524_/B sky130_fd_sc_hd__buf_2
XFILLER_54_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23731_ _24162_/CLK _23731_/D HRESETn VGND VGND VPWR VPWR _23731_/Q sky130_fd_sc_hd__dfrtp_4
X_20943_ _23938_/Q VGND VGND VPWR VPWR _20971_/A sky130_fd_sc_hd__buf_2
XANTENNA__12861__B2 _24459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25083__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18873__C _13461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23662_ _23661_/CLK _23662_/D HRESETn VGND VGND VPWR VPWR _23662_/Q sky130_fd_sc_hd__dfrtp_4
X_20874_ _14284_/Y _21590_/B _24772_/Q _21093_/B VGND VGND VPWR VPWR _20875_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14063__B1 _13398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25012__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22613_ _22360_/X _22593_/X _22597_/X _22604_/X _22612_/X VGND VGND VPWR VPWR _22613_/X
+ sky130_fd_sc_hd__o41a_4
XANTENNA__14475__A _14429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22676__A2 _22281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23593_ _23128_/CLK _23593_/D VGND VGND VPWR VPWR _13234_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16393__C _16041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22544_ _16430_/Y _22551_/A _14751_/Y _22225_/A VGND VGND VPWR VPWR _22544_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22692__A _24211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17786__A _17727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22475_ _12489_/A _22178_/X _24042_/Q _22260_/X VGND VGND VPWR VPWR _22476_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19829__B1 _19828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16690__A _22256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24214_ _23828_/CLK _16415_/X HRESETn VGND VGND VPWR VPWR _16413_/A sky130_fd_sc_hd__dfrtp_4
X_21426_ _22610_/A _21424_/X _21280_/X _21425_/X VGND VGND VPWR VPWR _21426_/X sky130_fd_sc_hd__o22a_4
X_25194_ _25194_/CLK _25194_/D HRESETn VGND VGND VPWR VPWR _25194_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21357_ _21357_/A VGND VGND VPWR VPWR _21357_/X sky130_fd_sc_hd__buf_2
XFILLER_135_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24145_ _24145_/CLK _16588_/X HRESETn VGND VGND VPWR VPWR _24145_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21458__D _21457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20308_ _14262_/Y _20296_/X _20287_/X _20307_/X VGND VGND VPWR VPWR _20309_/A sky130_fd_sc_hd__a211o_4
XFILLER_2_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12090_ _12172_/A _12088_/Y _25129_/Q _12089_/Y VGND VGND VPWR VPWR _12090_/X sky130_fd_sc_hd__a2bb2o_4
X_21288_ _13335_/X _21282_/X _22407_/A _21287_/X VGND VGND VPWR VPWR _21288_/X sky130_fd_sc_hd__o22a_4
XFILLER_1_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24076_ _24079_/CLK _16903_/X HRESETn VGND VGND VPWR VPWR _16784_/A sky130_fd_sc_hd__dfrtp_4
X_20239_ _20239_/A _20200_/A VGND VGND VPWR VPWR _20239_/X sky130_fd_sc_hd__and2_4
X_23027_ _21864_/X _23025_/Y _22530_/X _23026_/Y VGND VGND VPWR VPWR _23027_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19506__A _19859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18410__A _18484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23947__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14800_ _24683_/Q VGND VGND VPWR VPWR _15092_/A sky130_fd_sc_hd__inv_2
XFILLER_18_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15780_ _15748_/X _15763_/X _15494_/X _24445_/Q _15779_/X VGND VGND VPWR VPWR _24445_/D
+ sky130_fd_sc_hd__a32o_4
X_12992_ _12992_/A _12992_/B _12991_/Y VGND VGND VPWR VPWR _12992_/X sky130_fd_sc_hd__and3_4
X_24978_ _24980_/CLK _13380_/X HRESETn VGND VGND VPWR VPWR _24978_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22867__A _22931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14369__B _14369_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14731_ _24689_/Q VGND VGND VPWR VPWR _14844_/A sky130_fd_sc_hd__inv_2
XANTENNA__21771__A _21519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11943_ _22616_/A VGND VGND VPWR VPWR _22477_/B sky130_fd_sc_hd__buf_2
XFILLER_73_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23929_ _24735_/CLK _23929_/D HRESETn VGND VGND VPWR VPWR _23929_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22586__B _22435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17450_ _17449_/X VGND VGND VPWR VPWR _17452_/A sky130_fd_sc_hd__buf_2
XFILLER_75_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14662_ _14640_/X _14661_/X _15290_/A _14647_/X VGND VGND VPWR VPWR _14662_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__16159__A1_N _16157_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11874_ _11866_/X VGND VGND VPWR VPWR _11874_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14054__B1 _13668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16401_ _16401_/A VGND VGND VPWR VPWR _16426_/A sky130_fd_sc_hd__buf_2
X_13613_ _13613_/A _24616_/Q _11938_/A VGND VGND VPWR VPWR _13614_/A sky130_fd_sc_hd__or3_4
X_17381_ _17312_/C _17380_/X VGND VGND VPWR VPWR _17382_/D sky130_fd_sc_hd__or2_4
XFILLER_60_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14593_ _14592_/X VGND VGND VPWR VPWR _18719_/A sky130_fd_sc_hd__buf_2
XANTENNA__12604__B2 _24515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19120_ _18711_/X VGND VGND VPWR VPWR _19120_/X sky130_fd_sc_hd__buf_2
X_16332_ _24243_/Q VGND VGND VPWR VPWR _16332_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13544_ _20551_/B VGND VGND VPWR VPWR _20554_/B sky130_fd_sc_hd__inv_2
XFILLER_13_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20678__B2 _20602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19051_ _19051_/A VGND VGND VPWR VPWR _19051_/Y sky130_fd_sc_hd__inv_2
X_16263_ _14907_/Y _16257_/X _16261_/X _16262_/X VGND VGND VPWR VPWR _16263_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24735__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13475_ _13475_/A VGND VGND VPWR VPWR _13475_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_8_0_HCLK clkbuf_6_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18002_ _11688_/Y _17995_/X _16671_/X _17987_/A VGND VGND VPWR VPWR _23912_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20834__B _22228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12368__B1 _12498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15214_ _14969_/Y _15219_/A VGND VGND VPWR VPWR _15214_/Y sky130_fd_sc_hd__nand2_4
XFILLER_12_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12426_ _12399_/A VGND VGND VPWR VPWR _12442_/A sky130_fd_sc_hd__inv_2
X_16194_ _16193_/Y _16191_/X _15788_/X _16191_/X VGND VGND VPWR VPWR _24299_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22107__A _20961_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15145_ _15144_/X VGND VGND VPWR VPWR _15145_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15306__B1 HADDR[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12357_ _24472_/Q VGND VGND VPWR VPWR _12357_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15076_ _15067_/C _15079_/B VGND VGND VPWR VPWR _15077_/C sky130_fd_sc_hd__nand2_4
X_19953_ _19960_/A VGND VGND VPWR VPWR _19953_/X sky130_fd_sc_hd__buf_2
X_12288_ _12283_/B _12288_/B _12300_/C VGND VGND VPWR VPWR _25107_/D sky130_fd_sc_hd__and3_4
XFILLER_4_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14027_ _14025_/Y VGND VGND VPWR VPWR _14027_/X sky130_fd_sc_hd__buf_2
X_18904_ _18903_/Y _18900_/X _18880_/X _18900_/X VGND VGND VPWR VPWR _23525_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19884_ _19883_/X VGND VGND VPWR VPWR _19897_/A sky130_fd_sc_hd__inv_2
XANTENNA__16806__B1 _15830_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18835_ _23549_/Q VGND VGND VPWR VPWR _21947_/B sky130_fd_sc_hd__inv_2
XFILLER_45_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23688__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15978_ HWDATA[9] VGND VGND VPWR VPWR _15978_/X sky130_fd_sc_hd__buf_2
X_18766_ _17743_/B VGND VGND VPWR VPWR _18766_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23617__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22777__A _15271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14929_ _24273_/Q VGND VGND VPWR VPWR _14929_/Y sky130_fd_sc_hd__inv_2
X_17717_ _17717_/A VGND VGND VPWR VPWR _17727_/A sky130_fd_sc_hd__buf_2
XFILLER_64_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18697_ _18697_/A VGND VGND VPWR VPWR _18697_/X sky130_fd_sc_hd__buf_2
XFILLER_110_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12843__B2 _22463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17648_ _21336_/A _17648_/B VGND VGND VPWR VPWR _17648_/X sky130_fd_sc_hd__or2_4
X_17579_ _17578_/X VGND VGND VPWR VPWR _17580_/B sky130_fd_sc_hd__inv_2
XFILLER_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15793__B1 _15386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19318_ _13245_/B VGND VGND VPWR VPWR _19318_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20590_ _20590_/A _20590_/B VGND VGND VPWR VPWR _20590_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24476__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19249_ _21484_/B _19244_/X _11853_/X _19244_/X VGND VGND VPWR VPWR _23402_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22260_ _21434_/A VGND VGND VPWR VPWR _22260_/X sky130_fd_sc_hd__buf_2
XANTENNA__24405__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19287__B2 _19284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21211_ _21211_/A _21211_/B VGND VGND VPWR VPWR _21212_/C sky130_fd_sc_hd__or2_4
XFILLER_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21094__A1 _21275_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22191_ _11516_/B VGND VGND VPWR VPWR _22191_/X sky130_fd_sc_hd__buf_2
XANTENNA__21094__B2 _20863_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21142_ _21469_/A _21142_/B VGND VGND VPWR VPWR _21142_/X sky130_fd_sc_hd__or2_4
XFILLER_104_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20760__A _20759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21073_ _21073_/A _21113_/B VGND VGND VPWR VPWR _21073_/X sky130_fd_sc_hd__and2_4
XFILLER_115_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14520__B2 _14506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21397__A2 _21396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20024_ _23121_/Q VGND VGND VPWR VPWR _21460_/B sky130_fd_sc_hd__inv_2
X_24901_ _24902_/CLK _13913_/X HRESETn VGND VGND VPWR VPWR _13808_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_24_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21294__C _21432_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24832_ _24851_/CLK _14173_/Y HRESETn VGND VGND VPWR VPWR _18111_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22346__A1 _21529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_14_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24763_ _24968_/CLK _24763_/D HRESETn VGND VGND VPWR VPWR _13432_/A sky130_fd_sc_hd__dfrtp_4
X_21975_ _21972_/X _21973_/X _21974_/X _12075_/A _21187_/X VGND VGND VPWR VPWR _21975_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_27_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16685__A _16685_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20919__B _20866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23714_ _23744_/CLK _20506_/Y HRESETn VGND VGND VPWR VPWR _22656_/A sky130_fd_sc_hd__dfrtp_4
X_20926_ _20926_/A VGND VGND VPWR VPWR _20926_/X sky130_fd_sc_hd__buf_2
XPHY_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24694_ _24706_/CLK _15056_/Y HRESETn VGND VGND VPWR VPWR _14757_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_54_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15784__B1 _22385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23645_ _23796_/CLK sda_i_S4 HRESETn VGND VGND VPWR VPWR _23645_/Q sky130_fd_sc_hd__dfrtp_4
X_20857_ _24125_/Q _21297_/A VGND VGND VPWR VPWR _20857_/X sky130_fd_sc_hd__and2_4
XFILLER_74_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11590_ _16093_/A VGND VGND VPWR VPWR _11590_/X sky130_fd_sc_hd__buf_2
XPHY_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23576_ _23568_/CLK _23576_/D VGND VGND VPWR VPWR _18754_/A sky130_fd_sc_hd__dfxtp_4
X_20788_ _15653_/X VGND VGND VPWR VPWR _22953_/B sky130_fd_sc_hd__buf_2
XANTENNA__18722__B1 _18700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22527_ _22527_/A _22527_/B VGND VGND VPWR VPWR _22527_/X sky130_fd_sc_hd__and2_4
XFILLER_109_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_138_0_HCLK clkbuf_7_69_0_HCLK/X VGND VGND VPWR VPWR _23486_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13260_ _13122_/A _13258_/X _13259_/X VGND VGND VPWR VPWR _13260_/X sky130_fd_sc_hd__and3_4
XANTENNA__24146__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22458_ _22458_/A _22238_/X VGND VGND VPWR VPWR _22458_/X sky130_fd_sc_hd__or2_4
XFILLER_41_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12211_ _12185_/A _12209_/A VGND VGND VPWR VPWR _12211_/X sky130_fd_sc_hd__or2_4
X_21409_ _22501_/A _21408_/X _21036_/X _24548_/Q _11530_/X VGND VGND VPWR VPWR _21410_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21085__B2 _21425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13191_ _13113_/A _13180_/X _13191_/C VGND VGND VPWR VPWR _13191_/X sky130_fd_sc_hd__and3_4
X_25177_ _24847_/CLK _11825_/X HRESETn VGND VGND VPWR VPWR _11776_/B sky130_fd_sc_hd__dfrtp_4
X_22389_ _21042_/X _22388_/X _22197_/X _24408_/Q _20866_/X VGND VGND VPWR VPWR _22390_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_108_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12142_ _12171_/B _24567_/Q _12177_/A _12085_/Y VGND VGND VPWR VPWR _12142_/X sky130_fd_sc_hd__a2bb2o_4
X_24128_ _24104_/CLK _24128_/D HRESETn VGND VGND VPWR VPWR _24128_/Q sky130_fd_sc_hd__dfrtp_4
X_12073_ _25133_/Q VGND VGND VPWR VPWR _12073_/Y sky130_fd_sc_hd__inv_2
X_16950_ _16832_/Y _16953_/A VGND VGND VPWR VPWR _16950_/X sky130_fd_sc_hd__or2_4
X_24059_ _24064_/CLK _24059_/D HRESETn VGND VGND VPWR VPWR _24059_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_46_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15901_ _15899_/Y _15893_/X _15279_/X _15900_/X VGND VGND VPWR VPWR _15901_/X sky130_fd_sc_hd__a2bb2o_4
X_16881_ _16858_/A _16881_/B _16880_/X VGND VGND VPWR VPWR _16881_/X sky130_fd_sc_hd__or3_4
XANTENNA__20596__B1 _20583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13284__A _13316_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15832_ _24424_/Q VGND VGND VPWR VPWR _15832_/Y sky130_fd_sc_hd__inv_2
X_18620_ _18619_/X VGND VGND VPWR VPWR _18620_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23710__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15763_ _15740_/A VGND VGND VPWR VPWR _15763_/X sky130_fd_sc_hd__buf_2
X_18551_ _18551_/A _18551_/B VGND VGND VPWR VPWR _18552_/B sky130_fd_sc_hd__or2_4
XFILLER_79_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11516__B _11516_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12975_ _12974_/X VGND VGND VPWR VPWR _12976_/B sky130_fd_sc_hd__inv_2
XFILLER_131_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12825__B2 _21851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14714_ _14714_/A VGND VGND VPWR VPWR _14714_/Y sky130_fd_sc_hd__inv_2
X_17502_ _17481_/Y _17502_/B _17502_/C _17502_/D VGND VGND VPWR VPWR _17503_/B sky130_fd_sc_hd__or4_4
X_11926_ _11926_/A VGND VGND VPWR VPWR _21580_/A sky130_fd_sc_hd__inv_2
X_18482_ _18482_/A _18479_/B _18481_/X VGND VGND VPWR VPWR _18483_/A sky130_fd_sc_hd__or3_4
XFILLER_79_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15694_ _15693_/X _15689_/X _16100_/A _24478_/Q _15661_/A VGND VGND VPWR VPWR _15694_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24987__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16567__A2 _16276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17433_ _17433_/A VGND VGND VPWR VPWR _17433_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14645_ _23685_/D _14644_/X _20393_/A _23685_/D VGND VGND VPWR VPWR _24728_/D sky130_fd_sc_hd__a2bb2o_4
X_11857_ _19614_/A VGND VGND VPWR VPWR _11857_/X sky130_fd_sc_hd__buf_2
XANTENNA__24916__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11532__A _11532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17364_ _24001_/Q _17363_/Y VGND VGND VPWR VPWR _17364_/X sky130_fd_sc_hd__or2_4
X_14576_ _17717_/A VGND VGND VPWR VPWR _17729_/A sky130_fd_sc_hd__inv_2
XANTENNA__16651__A1_N _16649_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11788_ _11774_/Y _11785_/X _25185_/Q _11787_/X VGND VGND VPWR VPWR _25185_/D sky130_fd_sc_hd__o22a_4
XFILLER_14_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_34_0_HCLK clkbuf_7_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_69_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__21312__A2 _20931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16315_ _16312_/Y _16308_/X _16243_/X _16314_/X VGND VGND VPWR VPWR _16315_/X sky130_fd_sc_hd__a2bb2o_4
X_19103_ _17712_/B VGND VGND VPWR VPWR _19103_/Y sky130_fd_sc_hd__inv_2
X_13527_ _13525_/Y _13527_/B VGND VGND VPWR VPWR _13528_/A sky130_fd_sc_hd__and2_4
Xclkbuf_7_97_0_HCLK clkbuf_6_48_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_97_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17295_ _17291_/X _17295_/B _17293_/X _17294_/X VGND VGND VPWR VPWR _17296_/D sky130_fd_sc_hd__or4_4
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19034_ _19034_/A VGND VGND VPWR VPWR _19034_/Y sky130_fd_sc_hd__inv_2
X_16246_ HWDATA[27] VGND VGND VPWR VPWR _16246_/X sky130_fd_sc_hd__buf_2
X_13458_ _13471_/A _13458_/B VGND VGND VPWR VPWR _16035_/A sky130_fd_sc_hd__or2_4
XANTENNA__13002__A1 _12858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12409_ _12379_/Y _12409_/B _12409_/C _12505_/A VGND VGND VPWR VPWR _12409_/X sky130_fd_sc_hd__or4_4
XANTENNA__21076__B2 _15639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16177_ _16137_/A VGND VGND VPWR VPWR _16196_/A sky130_fd_sc_hd__buf_2
XFILLER_103_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13389_ _24976_/Q _20688_/B _13388_/X VGND VGND VPWR VPWR _13389_/X sky130_fd_sc_hd__a21o_4
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15128_ _15127_/X VGND VGND VPWR VPWR _24680_/D sky130_fd_sc_hd__inv_2
Xclkbuf_3_3_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__23869__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18229__C1 _18228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15059_ _15059_/A _15059_/B VGND VGND VPWR VPWR _15059_/X sky130_fd_sc_hd__or2_4
X_19936_ _23154_/Q VGND VGND VPWR VPWR _21502_/B sky130_fd_sc_hd__inv_2
XFILLER_130_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19867_ _21956_/B _19864_/X _19818_/X _19864_/X VGND VGND VPWR VPWR _23181_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18818_ _18816_/Y _18814_/X _18817_/X _18814_/X VGND VGND VPWR VPWR _18818_/X sky130_fd_sc_hd__a2bb2o_4
X_19798_ _19797_/Y _19793_/X _19506_/X _19780_/Y VGND VGND VPWR VPWR _23207_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22328__A1 _16445_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16604__A1_N _14831_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22938__C _22931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18749_ _17864_/B VGND VGND VPWR VPWR _18749_/Y sky130_fd_sc_hd__inv_2
X_21760_ _14443_/B VGND VGND VPWR VPWR _21760_/X sky130_fd_sc_hd__buf_2
XFILLER_37_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20711_ _20710_/A _13923_/B _20710_/C VGND VGND VPWR VPWR _20711_/X sky130_fd_sc_hd__or3_4
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15766__B1 _15765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24657__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21691_ _19268_/Y _21638_/X _19220_/Y _21795_/B VGND VGND VPWR VPWR _21691_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12538__A _12322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23430_ _23596_/CLK _19171_/X VGND VGND VPWR VPWR _23430_/Q sky130_fd_sc_hd__dfxtp_4
X_20642_ _20642_/A VGND VGND VPWR VPWR _20642_/Y sky130_fd_sc_hd__inv_2
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20755__A _13614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21303__A2 _20751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20573_ _20573_/A VGND VGND VPWR VPWR _23731_/D sky130_fd_sc_hd__inv_2
XFILLER_108_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15849__A _15849_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23361_ _25002_/CLK _23361_/D VGND VGND VPWR VPWR _19362_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__14959__A2_N _24281_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25100_ _23716_/CLK _12429_/Y HRESETn VGND VGND VPWR VPWR _12391_/A sky130_fd_sc_hd__dfrtp_4
X_22312_ _22312_/A _22312_/B VGND VGND VPWR VPWR _22312_/Y sky130_fd_sc_hd__nor2_4
XFILLER_30_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23292_ _23292_/CLK _23292_/D VGND VGND VPWR VPWR _23292_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_121_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25031_ _24451_/CLK _12914_/Y HRESETn VGND VGND VPWR VPWR _22854_/A sky130_fd_sc_hd__dfrtp_4
X_22243_ _22243_/A _20787_/B VGND VGND VPWR VPWR _22243_/X sky130_fd_sc_hd__or2_4
XANTENNA__14741__A1 _24711_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14741__B2 _14740_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22174_ _16700_/X _22637_/A _20590_/A _22173_/X VGND VGND VPWR VPWR _22174_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21125_ _13357_/X _21124_/X _21432_/C _24396_/Q _21285_/B VGND VGND VPWR VPWR _21126_/C
+ sky130_fd_sc_hd__a32o_4
XFILLER_78_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24805__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24868__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21056_ _21034_/Y VGND VGND VPWR VPWR _21432_/C sky130_fd_sc_hd__buf_2
XFILLER_87_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20007_ _20007_/A VGND VGND VPWR VPWR _20007_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24815_ _23774_/CLK _14229_/X HRESETn VGND VGND VPWR VPWR _14223_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__12807__A1 _22133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17304__A _17303_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12760_ _12737_/A _12737_/B _12758_/B _12674_/X VGND VGND VPWR VPWR _12761_/A sky130_fd_sc_hd__a211o_4
XPHY_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24746_ _25052_/CLK _24746_/D HRESETn VGND VGND VPWR VPWR _24746_/Q sky130_fd_sc_hd__dfrtp_4
X_21958_ _14524_/A _21956_/X _21957_/X VGND VGND VPWR VPWR _21958_/X sky130_fd_sc_hd__and3_4
XANTENNA__23025__B _23025_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11710_/X VGND VGND VPWR VPWR _11711_/X sky130_fd_sc_hd__buf_2
XFILLER_37_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ _13358_/X VGND VGND VPWR VPWR _20909_/X sky130_fd_sc_hd__buf_2
XANTENNA__24398__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12637_/X _12691_/B _12690_/Y VGND VGND VPWR VPWR _25061_/D sky130_fd_sc_hd__and3_4
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24677_ _24676_/CLK _24677_/D HRESETn VGND VGND VPWR VPWR _24677_/Q sky130_fd_sc_hd__dfrtp_4
X_21889_ _21887_/Y _13335_/X _22407_/A _21888_/X VGND VGND VPWR VPWR _21890_/B sky130_fd_sc_hd__o22a_4
XANTENNA__12448__A _12448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14430_/A VGND VGND VPWR VPWR _21403_/A sky130_fd_sc_hd__inv_2
XPHY_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _13644_/A VGND VGND VPWR VPWR _11643_/A sky130_fd_sc_hd__buf_2
XANTENNA__24327__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23628_ _23624_/CLK _20709_/A HRESETn VGND VGND VPWR VPWR _20710_/C sky130_fd_sc_hd__dfstp_4
XFILLER_39_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ _13840_/Y _14361_/B _14361_/C _14360_/X VGND VGND VPWR VPWR _14362_/A sky130_fd_sc_hd__or4_4
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11573_ HWDATA[17] VGND VGND VPWR VPWR _11573_/X sky130_fd_sc_hd__buf_2
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23559_ _23586_/CLK _23559_/D VGND VGND VPWR VPWR _17957_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16100_ _16100_/A VGND VGND VPWR VPWR _16100_/X sky130_fd_sc_hd__buf_2
XFILLER_122_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ _13092_/A _19391_/A VGND VGND VPWR VPWR _13312_/X sky130_fd_sc_hd__or2_4
XFILLER_11_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17080_ _17080_/A _17079_/Y VGND VGND VPWR VPWR _17080_/X sky130_fd_sc_hd__or2_4
X_14292_ _24789_/Q VGND VGND VPWR VPWR _14292_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16182__B1 _16087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22880__A _24217_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16031_ _17702_/A _16030_/Y _17702_/A _16030_/Y VGND VGND VPWR VPWR _16032_/A sky130_fd_sc_hd__a2bb2o_4
X_13243_ _13090_/X _13243_/B _13243_/C VGND VGND VPWR VPWR _13243_/X sky130_fd_sc_hd__and3_4
XANTENNA__13279__A _13073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21496__A _13337_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20805__B2 _20802_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13174_ _13136_/A _23371_/Q VGND VGND VPWR VPWR _13174_/X sky130_fd_sc_hd__or2_4
XANTENNA__23962__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12125_ _24550_/Q VGND VGND VPWR VPWR _12125_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22007__B1 _22005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15494__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17982_ _17982_/A VGND VGND VPWR VPWR _17982_/X sky130_fd_sc_hd__buf_2
XFILLER_2_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25115__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19721_ _11842_/A VGND VGND VPWR VPWR _19721_/X sky130_fd_sc_hd__buf_2
X_12056_ _12055_/X VGND VGND VPWR VPWR _12056_/Y sky130_fd_sc_hd__inv_2
X_16933_ _16927_/A _16936_/B VGND VGND VPWR VPWR _16934_/C sky130_fd_sc_hd__nand2_4
XFILLER_77_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19652_ _19646_/Y VGND VGND VPWR VPWR _19652_/X sky130_fd_sc_hd__buf_2
X_16864_ _16866_/B VGND VGND VPWR VPWR _16864_/Y sky130_fd_sc_hd__inv_2
X_18603_ _18587_/X _18592_/X _18603_/C _18602_/X VGND VGND VPWR VPWR _18603_/X sky130_fd_sc_hd__or4_4
XFILLER_37_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15815_ _15814_/X VGND VGND VPWR VPWR _15815_/Y sky130_fd_sc_hd__inv_2
X_16795_ _15870_/Y _16824_/A _15870_/Y _16824_/A VGND VGND VPWR VPWR _16795_/X sky130_fd_sc_hd__a2bb2o_4
X_19583_ _19583_/A VGND VGND VPWR VPWR _21674_/B sky130_fd_sc_hd__inv_2
XFILLER_24_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15996__B1 _15282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22120__A _22438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15746_ _15746_/A VGND VGND VPWR VPWR _15746_/X sky130_fd_sc_hd__buf_2
X_18534_ _18534_/A VGND VGND VPWR VPWR _23823_/D sky130_fd_sc_hd__inv_2
X_12958_ _12880_/A _12955_/X VGND VGND VPWR VPWR _12958_/X sky130_fd_sc_hd__or2_4
XFILLER_18_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11909_ _23789_/Q _11905_/X VGND VGND VPWR VPWR _11909_/X sky130_fd_sc_hd__and2_4
XANTENNA__13461__B _13460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24750__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15677_ _15666_/A VGND VGND VPWR VPWR _15677_/X sky130_fd_sc_hd__buf_2
X_18465_ _18438_/B _18445_/X _18438_/A VGND VGND VPWR VPWR _18465_/X sky130_fd_sc_hd__o21a_4
X_12889_ _23013_/A _12888_/Y VGND VGND VPWR VPWR _12889_/X sky130_fd_sc_hd__or2_4
X_14628_ _24726_/Q _14627_/X _24727_/Q VGND VGND VPWR VPWR _14628_/X sky130_fd_sc_hd__or3_4
X_17416_ _17319_/Y _17419_/B _17336_/X VGND VGND VPWR VPWR _17416_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24068__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18396_ _16464_/Y _18419_/A _24218_/Q _18452_/C VGND VGND VPWR VPWR _18401_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17347_ _17347_/A VGND VGND VPWR VPWR _24006_/D sky130_fd_sc_hd__inv_2
X_14559_ _14563_/A _14558_/X VGND VGND VPWR VPWR _14560_/A sky130_fd_sc_hd__and2_4
XFILLER_18_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18162__A1 _16078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14971__B2 _24258_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17278_ _11587_/Y _17315_/A _11587_/Y _17315_/A VGND VGND VPWR VPWR _17278_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16173__B1 _15775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_121_0_HCLK clkbuf_7_60_0_HCLK/X VGND VGND VPWR VPWR _23845_/CLK sky130_fd_sc_hd__clkbuf_1
X_16229_ _11949_/Y _14195_/B _14195_/C _16038_/D VGND VGND VPWR VPWR _20856_/A sky130_fd_sc_hd__or4_4
X_19017_ _23484_/Q VGND VGND VPWR VPWR _21769_/B sky130_fd_sc_hd__inv_2
XFILLER_127_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_184_0_HCLK clkbuf_7_92_0_HCLK/X VGND VGND VPWR VPWR _25123_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22797__A1 _15821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16476__A1 _15619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12821__A _12811_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23632__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22014__B _22014_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19919_ _19917_/Y _19918_/X _19832_/X _19918_/X VGND VGND VPWR VPWR _19919_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19414__B2 _19396_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20805__A1_N _20802_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19604__A _19613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22930_ _24250_/Q _16134_/X _22858_/X _22929_/X VGND VGND VPWR VPWR _22930_/X sky130_fd_sc_hd__a211o_4
XFILLER_99_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24838__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22861_ _14859_/A _15919_/X _22858_/X _22860_/X VGND VGND VPWR VPWR _22862_/C sky130_fd_sc_hd__a211o_4
XANTENNA__19178__B1 _19109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24600_ _24606_/CLK _15364_/X HRESETn VGND VGND VPWR VPWR _15363_/A sky130_fd_sc_hd__dfrtp_4
X_21812_ _20966_/A _21812_/B VGND VGND VPWR VPWR _21812_/X sky130_fd_sc_hd__or2_4
XANTENNA__17124__A _17053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22792_ _14850_/Y _21043_/X _14913_/Y _22154_/B VGND VGND VPWR VPWR _22792_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18925__B1 _18880_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24531_ _25005_/CLK _24531_/D HRESETn VGND VGND VPWR VPWR _12579_/A sky130_fd_sc_hd__dfrtp_4
X_21743_ _21739_/X _21740_/X _21741_/X _21742_/X VGND VGND VPWR VPWR _21743_/X sky130_fd_sc_hd__or4_4
XANTENNA__15739__B1 _24462_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24491__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24420__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24462_ _24944_/CLK _24462_/D HRESETn VGND VGND VPWR VPWR _24462_/Q sky130_fd_sc_hd__dfrtp_4
X_21674_ _21205_/A _21674_/B VGND VGND VPWR VPWR _21674_/X sky130_fd_sc_hd__or2_4
XANTENNA__20485__A _13509_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21288__A1 _13335_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23413_ _23085_/CLK _23413_/D VGND VGND VPWR VPWR _21876_/A sky130_fd_sc_hd__dfxtp_4
X_20625_ _20621_/X _20623_/Y _24173_/Q _20624_/X VGND VGND VPWR VPWR _23742_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24393_ _24071_/CLK _15914_/X HRESETn VGND VGND VPWR VPWR _24393_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17497__C _16692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23344_ _23336_/CLK _19412_/X VGND VGND VPWR VPWR _19411_/A sky130_fd_sc_hd__dfxtp_4
X_20556_ _20647_/A VGND VGND VPWR VPWR _20556_/X sky130_fd_sc_hd__buf_2
XFILLER_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_80_0_HCLK clkbuf_6_40_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_80_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15506__A3 _15505_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16703__A2 _22782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13099__A _13316_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23275_ _23353_/CLK _19608_/X VGND VGND VPWR VPWR _19606_/A sky130_fd_sc_hd__dfxtp_4
X_20487_ _13509_/A _20481_/X _20495_/B VGND VGND VPWR VPWR _20487_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_106_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22788__B2 _21069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25014_ _24435_/CLK _12986_/X HRESETn VGND VGND VPWR VPWR _22203_/A sky130_fd_sc_hd__dfrtp_4
X_22226_ _22226_/A VGND VGND VPWR VPWR _22226_/X sky130_fd_sc_hd__buf_2
XFILLER_105_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22252__A3 _22251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12825__A1_N _12951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22205__A _21175_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22157_ _22157_/A VGND VGND VPWR VPWR _22168_/A sky130_fd_sc_hd__inv_2
XFILLER_65_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21108_ _21104_/X _21105_/X _21107_/X VGND VGND VPWR VPWR _21108_/X sky130_fd_sc_hd__o21a_4
X_22088_ _20946_/X _19594_/Y VGND VGND VPWR VPWR _22088_/X sky130_fd_sc_hd__or2_4
XFILLER_134_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20021__A2_N _20015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17416__B1 _17336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13930_ _24892_/Q _13930_/B _13939_/A VGND VGND VPWR VPWR _13930_/X sky130_fd_sc_hd__or3_4
XFILLER_102_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21039_ _11516_/B VGND VGND VPWR VPWR _22637_/A sky130_fd_sc_hd__buf_2
XFILLER_75_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23681__D scl_i_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22960__B2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13861_ _13861_/A _13812_/X _13872_/A _13851_/X VGND VGND VPWR VPWR _13862_/A sky130_fd_sc_hd__or4_4
XANTENNA__24579__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15600_ HWDATA[23] VGND VGND VPWR VPWR _15600_/X sky130_fd_sc_hd__buf_2
X_12812_ _12812_/A VGND VGND VPWR VPWR _12812_/Y sky130_fd_sc_hd__inv_2
X_16580_ _14850_/Y _16576_/X _16251_/X _16576_/X VGND VGND VPWR VPWR _24149_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24508__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13792_ _13744_/X _13792_/B _13792_/C VGND VGND VPWR VPWR _13793_/B sky130_fd_sc_hd__or3_4
XFILLER_28_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15531_ _16302_/A _15531_/B VGND VGND VPWR VPWR _15531_/X sky130_fd_sc_hd__or2_4
X_12743_ _12648_/Y _12742_/X VGND VGND VPWR VPWR _12747_/B sky130_fd_sc_hd__or2_4
X_24729_ _23661_/CLK _14642_/X HRESETn VGND VGND VPWR VPWR _24729_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_76_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18250_ _18242_/B _18257_/B VGND VGND VPWR VPWR _18250_/X sky130_fd_sc_hd__or2_4
X_15462_ _13357_/X VGND VGND VPWR VPWR _15463_/A sky130_fd_sc_hd__buf_2
XANTENNA__24161__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12674_ _13007_/B VGND VGND VPWR VPWR _12674_/X sky130_fd_sc_hd__buf_2
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _24018_/Q VGND VGND VPWR VPWR _17201_/Y sky130_fd_sc_hd__inv_2
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14380_/X _14411_/Y _14412_/X _14403_/X _13413_/A VGND VGND VPWR VPWR _14413_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _11625_/A VGND VGND VPWR VPWR _13632_/A sky130_fd_sc_hd__buf_2
X_18181_ _23865_/Q VGND VGND VPWR VPWR _18207_/B sky130_fd_sc_hd__inv_2
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ _16376_/A VGND VGND VPWR VPWR _15393_/X sky130_fd_sc_hd__buf_2
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17132_ _17132_/A _17035_/C VGND VGND VPWR VPWR _17133_/B sky130_fd_sc_hd__or2_4
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14344_ _24773_/Q _14325_/A _24772_/Q _14319_/X VGND VGND VPWR VPWR _14344_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21597__A1_N _12972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11556_ _11554_/Y _11551_/X _11555_/X _11551_/X VGND VGND VPWR VPWR _25213_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17063_ _17022_/A _17063_/B VGND VGND VPWR VPWR _17064_/C sky130_fd_sc_hd__or2_4
XFILLER_6_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14275_ _24796_/Q VGND VGND VPWR VPWR _14275_/Y sky130_fd_sc_hd__inv_2
X_16014_ _16014_/A _16014_/B _16014_/C VGND VGND VPWR VPWR _16014_/X sky130_fd_sc_hd__and3_4
XFILLER_100_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13226_ _11732_/B _13226_/B VGND VGND VPWR VPWR _13226_/X sky130_fd_sc_hd__or2_4
X_13157_ _13120_/X _13157_/B VGND VGND VPWR VPWR _13157_/X sky130_fd_sc_hd__or2_4
XFILLER_88_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12108_ _24574_/Q VGND VGND VPWR VPWR _12108_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13456__B _14369_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13088_ _13011_/X _13073_/X _13088_/C VGND VGND VPWR VPWR _13088_/X sky130_fd_sc_hd__and3_4
X_17965_ _17716_/X _17963_/X _17965_/C VGND VGND VPWR VPWR _17969_/B sky130_fd_sc_hd__and3_4
X_19704_ _19703_/Y _19701_/X _19617_/X _19701_/X VGND VGND VPWR VPWR _19704_/X sky130_fd_sc_hd__a2bb2o_4
X_12039_ _12039_/A _12035_/X VGND VGND VPWR VPWR _12041_/A sky130_fd_sc_hd__and2_4
X_16916_ _16916_/A _16916_/B VGND VGND VPWR VPWR _16917_/C sky130_fd_sc_hd__or2_4
XFILLER_78_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19424__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17896_ _17928_/A _23577_/Q VGND VGND VPWR VPWR _17897_/C sky130_fd_sc_hd__or2_4
XFILLER_77_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19635_ _23265_/Q VGND VGND VPWR VPWR _21335_/B sky130_fd_sc_hd__inv_2
X_16847_ _16867_/A _16845_/X _16846_/Y VGND VGND VPWR VPWR _24090_/D sky130_fd_sc_hd__and3_4
XANTENNA__15969__B1 _11590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24931__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14568__A _17732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13472__A _13461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24249__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19566_ _23289_/Q VGND VGND VPWR VPWR _21344_/B sky130_fd_sc_hd__inv_2
XFILLER_53_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16778_ _24061_/Q VGND VGND VPWR VPWR _16778_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_5_23_0_HCLK_A clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14287__B _18633_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18517_ _18517_/A _18517_/B VGND VGND VPWR VPWR _18519_/B sky130_fd_sc_hd__or2_4
XFILLER_20_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15729_ _15729_/A VGND VGND VPWR VPWR _15729_/X sky130_fd_sc_hd__buf_2
X_19497_ _21654_/B _19494_/X _19452_/X _19494_/X VGND VGND VPWR VPWR _19497_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12088__A _12088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18448_ _18448_/A VGND VGND VPWR VPWR _18475_/A sky130_fd_sc_hd__inv_2
XFILLER_21_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19299__A2_N _19296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22467__B1 _24410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18379_ _18503_/A VGND VGND VPWR VPWR _18495_/B sky130_fd_sc_hd__inv_2
XANTENNA__19332__B1 _19308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20410_ _20410_/A VGND VGND VPWR VPWR _23688_/D sky130_fd_sc_hd__inv_2
X_21390_ _21235_/A _19792_/Y VGND VGND VPWR VPWR _21390_/X sky130_fd_sc_hd__or2_4
XANTENNA__16146__B1 _15753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12624__A2_N _24505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23884__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20341_ _20198_/X _20234_/X VGND VGND VPWR VPWR _23652_/D sky130_fd_sc_hd__and2_4
XANTENNA__21848__B _21848_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23813__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25037__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20272_ _18622_/X VGND VGND VPWR VPWR _20296_/A sky130_fd_sc_hd__inv_2
X_23060_ _20738_/X VGND VGND VPWR VPWR IRQ[8] sky130_fd_sc_hd__buf_2
XFILLER_108_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22011_ _22011_/A VGND VGND VPWR VPWR _22011_/X sky130_fd_sc_hd__buf_2
XFILLER_103_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13380__B1 _11981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21864__A _22279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15862__A _15862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21583__B _21582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23962_ _23957_/CLK _23962_/D HRESETn VGND VGND VPWR VPWR _23962_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22913_ _22913_/A _22015_/X VGND VGND VPWR VPWR _22913_/X sky130_fd_sc_hd__or2_4
XANTENNA__24672__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23893_ _23990_/CLK _23893_/D HRESETn VGND VGND VPWR VPWR _23893_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_83_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24601__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22844_ _24455_/Q _22015_/X VGND VGND VPWR VPWR _22844_/X sky130_fd_sc_hd__or2_4
XFILLER_73_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22775_ _22775_/A _22756_/X _22661_/C _22775_/D VGND VGND VPWR VPWR HRDATA[23] sky130_fd_sc_hd__or4_4
XANTENNA__16693__A _16693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18374__A1 _16450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24514_ _24483_/CLK _24514_/D HRESETn VGND VGND VPWR VPWR _24514_/Q sky130_fd_sc_hd__dfrtp_4
X_21726_ _21724_/X _21725_/X _11532_/A VGND VGND VPWR VPWR _21726_/X sky130_fd_sc_hd__o21a_4
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21104__A _21104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24445_ _24445_/CLK _24445_/D HRESETn VGND VGND VPWR VPWR _24445_/Q sky130_fd_sc_hd__dfrtp_4
X_21657_ _21657_/A _21657_/B VGND VGND VPWR VPWR _21660_/B sky130_fd_sc_hd__or2_4
XFILLER_138_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11630__A _11630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20608_ _20598_/X _20607_/X _16527_/A _20603_/X VGND VGND VPWR VPWR _20608_/X sky130_fd_sc_hd__a2bb2o_4
X_12390_ _12389_/X _24470_/Q _21104_/A _12356_/Y VGND VGND VPWR VPWR _12390_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14760__A2_N _24107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24376_ _24372_/CLK _15962_/X HRESETn VGND VGND VPWR VPWR _22521_/A sky130_fd_sc_hd__dfrtp_4
X_21588_ _11952_/X _21582_/X VGND VGND VPWR VPWR _21881_/A sky130_fd_sc_hd__or2_4
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23327_ _24740_/CLK _19465_/X VGND VGND VPWR VPWR _19464_/A sky130_fd_sc_hd__dfxtp_4
X_20539_ _20542_/B _13514_/X _20538_/Y VGND VGND VPWR VPWR _20539_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__21758__B _23034_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14060_ _14048_/A VGND VGND VPWR VPWR _14060_/X sky130_fd_sc_hd__buf_2
X_23258_ _23258_/CLK _23258_/D VGND VGND VPWR VPWR _19656_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_106_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13011_ _23893_/Q VGND VGND VPWR VPWR _13011_/X sky130_fd_sc_hd__buf_2
XANTENNA__13371__B1 _11620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22209_ _22206_/X _22208_/X _11532_/X VGND VGND VPWR VPWR _22209_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17637__B1 _17636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22630__B1 _24564_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23189_ _23179_/CLK _23189_/D VGND VGND VPWR VPWR _23189_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_24_0_HCLK clkbuf_7_12_0_HCLK/X VGND VGND VPWR VPWR _24750_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_87_0_HCLK clkbuf_8_87_0_HCLK/A VGND VGND VPWR VPWR _24902_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_95_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15663__A2 _15647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15772__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14962_ _24672_/Q _14960_/Y _15161_/A _24275_/Q VGND VGND VPWR VPWR _14962_/X sky130_fd_sc_hd__a2bb2o_4
X_17750_ _17935_/A _17750_/B VGND VGND VPWR VPWR _17750_/X sky130_fd_sc_hd__or2_4
XFILLER_75_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16701_ _15981_/A _16699_/A _15981_/Y _16700_/X VGND VGND VPWR VPWR _16707_/B sky130_fd_sc_hd__o22a_4
X_13913_ _23693_/Q _13905_/A _13900_/X _13808_/X _13911_/X VGND VGND VPWR VPWR _13913_/X
+ sky130_fd_sc_hd__a32o_4
X_14893_ _14884_/X _14886_/X _14889_/X _14893_/D VGND VGND VPWR VPWR _14893_/X sky130_fd_sc_hd__or4_4
X_17681_ _17697_/A _17681_/B VGND VGND VPWR VPWR _17681_/X sky130_fd_sc_hd__or2_4
XFILLER_63_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19420_ _23341_/Q VGND VGND VPWR VPWR _19420_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13292__A _11751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13844_ _13829_/X VGND VGND VPWR VPWR _13844_/Y sky130_fd_sc_hd__inv_2
X_16632_ _16632_/A VGND VGND VPWR VPWR _16632_/X sky130_fd_sc_hd__buf_2
XFILLER_75_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24342__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19351_ _19347_/Y _19350_/X _19329_/X _19350_/X VGND VGND VPWR VPWR _19351_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13775_ _13762_/D VGND VGND VPWR VPWR _13775_/Y sky130_fd_sc_hd__inv_2
X_16563_ _20863_/A VGND VGND VPWR VPWR _23008_/B sky130_fd_sc_hd__buf_2
XANTENNA__22697__B1 _21562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18302_ _18216_/A _18321_/A VGND VGND VPWR VPWR _18302_/X sky130_fd_sc_hd__or2_4
X_12726_ _12636_/X VGND VGND VPWR VPWR _12749_/A sky130_fd_sc_hd__buf_2
X_15514_ _15470_/Y VGND VGND VPWR VPWR _15514_/X sky130_fd_sc_hd__buf_2
X_16494_ _16492_/Y _16493_/X _15479_/X _16493_/X VGND VGND VPWR VPWR _16494_/X sky130_fd_sc_hd__a2bb2o_4
X_19282_ _18018_/X _19282_/B _18031_/C VGND VGND VPWR VPWR _19283_/A sky130_fd_sc_hd__or3_4
XFILLER_31_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15445_ _14433_/X _15441_/B _15449_/B VGND VGND VPWR VPWR _15445_/Y sky130_fd_sc_hd__o21ai_4
X_18233_ _18232_/X VGND VGND VPWR VPWR _18234_/B sky130_fd_sc_hd__inv_2
X_12657_ _12657_/A _12727_/A _12641_/X _12663_/A VGND VGND VPWR VPWR _12657_/X sky130_fd_sc_hd__or4_4
XFILLER_128_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11540__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11608_ _11606_/Y _11599_/X _11607_/X _11599_/X VGND VGND VPWR VPWR _25198_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15376_ _24595_/Q VGND VGND VPWR VPWR _22323_/A sky130_fd_sc_hd__inv_2
X_18164_ _18164_/A _18164_/B _18154_/X _18163_/X VGND VGND VPWR VPWR _18164_/X sky130_fd_sc_hd__or4_4
XANTENNA__21949__A _21374_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12588_ _12588_/A VGND VGND VPWR VPWR _12588_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21121__B1 _21179_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20853__A _11503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14327_ _14315_/C VGND VGND VPWR VPWR _14327_/X sky130_fd_sc_hd__buf_2
X_17115_ _17115_/A VGND VGND VPWR VPWR _24043_/D sky130_fd_sc_hd__inv_2
X_11539_ _25217_/Q VGND VGND VPWR VPWR _11539_/Y sky130_fd_sc_hd__inv_2
X_18095_ _11767_/X _18095_/B VGND VGND VPWR VPWR _18095_/X sky130_fd_sc_hd__or2_4
XFILLER_8_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25130__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17046_ _17023_/Y _17045_/X VGND VGND VPWR VPWR _17046_/X sky130_fd_sc_hd__or2_4
X_14258_ _14257_/Y _14253_/X _14221_/X _14253_/X VGND VGND VPWR VPWR _14258_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13209_ _13136_/A _23370_/Q VGND VGND VPWR VPWR _13209_/X sky130_fd_sc_hd__or2_4
XFILLER_124_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14189_ _14174_/Y _14188_/X _25150_/Q _14180_/X VGND VGND VPWR VPWR _24826_/D sky130_fd_sc_hd__o22a_4
XFILLER_135_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18997_ _21763_/B _18991_/X _15550_/X _18996_/X VGND VGND VPWR VPWR _18997_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17948_ _17916_/A _17948_/B VGND VGND VPWR VPWR _17948_/X sky130_fd_sc_hd__or2_4
XFILLER_66_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17879_ _17879_/A _17877_/X _17879_/C VGND VGND VPWR VPWR _17883_/B sky130_fd_sc_hd__and3_4
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19618_ _21146_/B _19613_/X _19617_/X _19613_/X VGND VGND VPWR VPWR _23272_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24083__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20890_ _20885_/X _20888_/X _11954_/A _20889_/X VGND VGND VPWR VPWR _20890_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24012__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19549_ _19548_/Y _19546_/X _11860_/X _19546_/X VGND VGND VPWR VPWR _19549_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16367__B1 _15982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22560_ _24306_/Q _22957_/B VGND VGND VPWR VPWR _22560_/X sky130_fd_sc_hd__and2_4
X_21511_ _21507_/X _21510_/X _21242_/X VGND VGND VPWR VPWR _21511_/X sky130_fd_sc_hd__o21a_4
X_22491_ _23742_/Q _22173_/X _13509_/A _22170_/X VGND VGND VPWR VPWR _22491_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__14917__B2 _14916_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25218__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24230_ _23840_/CLK _24230_/D HRESETn VGND VGND VPWR VPWR _16366_/A sky130_fd_sc_hd__dfrtp_4
X_21442_ _21441_/X VGND VGND VPWR VPWR _21457_/B sky130_fd_sc_hd__inv_2
XFILLER_119_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21112__B1 _22279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14238__A1_N _14234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20763__A _11940_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11600__B1 _11598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15857__A _24415_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24161_ _24161_/CLK _24161_/D HRESETn VGND VGND VPWR VPWR _16548_/A sky130_fd_sc_hd__dfrtp_4
X_21373_ _21369_/X _21372_/X _21231_/X VGND VGND VPWR VPWR _21373_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19329__A _18763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23112_ _23112_/CLK _20049_/X VGND VGND VPWR VPWR _20047_/A sky130_fd_sc_hd__dfxtp_4
X_20324_ _23640_/Q _18617_/X _20323_/Y _20296_/A VGND VGND VPWR VPWR _20324_/X sky130_fd_sc_hd__a211o_4
XFILLER_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24092_ _23990_/CLK _24092_/D HRESETn VGND VGND VPWR VPWR _13461_/C sky130_fd_sc_hd__dfrtp_4
XANTENNA__21415__A1 _15322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12156__B2 _24549_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23043_ _22263_/X _15920_/A HWDATA[31] _25221_/Q _11537_/X VGND VGND VPWR VPWR _23043_/X
+ sky130_fd_sc_hd__a32o_4
X_20255_ _20254_/X VGND VGND VPWR VPWR _20255_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_240_0_HCLK clkbuf_8_241_0_HCLK/A VGND VGND VPWR VPWR _24140_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__11903__A1 _22006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21594__A _17027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20186_ _23691_/Q _20251_/B _20179_/X _20185_/Y VGND VGND VPWR VPWR _20186_/X sky130_fd_sc_hd__a211o_4
XFILLER_27_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24853__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24994_ _24841_/CLK _24994_/D HRESETn VGND VGND VPWR VPWR _13332_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22202__B _22438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23945_ _23972_/CLK _23945_/D HRESETn VGND VGND VPWR VPWR _23945_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14806__A1_N _14703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11625__A _11625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11890_ _11890_/A VGND VGND VPWR VPWR _11890_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23876_ _24641_/CLK _23876_/D HRESETn VGND VGND VPWR VPWR _23876_/Q sky130_fd_sc_hd__dfrtp_4
X_22827_ _12451_/A _22606_/X _17080_/A _22652_/X VGND VGND VPWR VPWR _22830_/B sky130_fd_sc_hd__a2bb2o_4
X_13560_ _13591_/A _13559_/X VGND VGND VPWR VPWR _13561_/B sky130_fd_sc_hd__or2_4
XANTENNA__19744__A2_N _19738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22758_ _22195_/X _22757_/X _22629_/X _24568_/Q _22198_/X VGND VGND VPWR VPWR _22759_/B
+ sky130_fd_sc_hd__a32o_4
X_12511_ _12345_/X _12328_/Y _12407_/B _12511_/D VGND VGND VPWR VPWR _12511_/X sky130_fd_sc_hd__or4_4
XFILLER_129_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21709_ _21434_/A VGND VGND VPWR VPWR _22968_/A sky130_fd_sc_hd__buf_2
X_13491_ _20883_/A _14106_/B VGND VGND VPWR VPWR _13492_/A sky130_fd_sc_hd__or2_4
XANTENNA__23735__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22689_ _14900_/A _22616_/X _22338_/X VGND VGND VPWR VPWR _22689_/X sky130_fd_sc_hd__o21a_4
X_15230_ _24651_/Q _15230_/B VGND VGND VPWR VPWR _15231_/B sky130_fd_sc_hd__or2_4
X_12442_ _12442_/A VGND VGND VPWR VPWR _12444_/A sky130_fd_sc_hd__buf_2
XFILLER_90_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24428_ _23442_/CLK _15816_/X HRESETn VGND VGND VPWR VPWR _15807_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_12_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15161_ _15161_/A _15161_/B VGND VGND VPWR VPWR _15162_/A sky130_fd_sc_hd__or2_4
XANTENNA__12395__B2 _24470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12373_ _12373_/A VGND VGND VPWR VPWR _12411_/A sky130_fd_sc_hd__inv_2
X_24359_ _23353_/CLK _16015_/X HRESETn VGND VGND VPWR VPWR _24359_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_50_0_HCLK clkbuf_6_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_50_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14112_ _14111_/X VGND VGND VPWR VPWR _14112_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15092_ _15092_/A _15085_/X VGND VGND VPWR VPWR _15093_/C sky130_fd_sc_hd__nand2_4
XFILLER_4_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14043_ _20405_/A VGND VGND VPWR VPWR _14043_/Y sky130_fd_sc_hd__inv_2
X_18920_ _18920_/A _19144_/B _19100_/A VGND VGND VPWR VPWR _18920_/X sky130_fd_sc_hd__or3_4
XANTENNA__21406__A1 _21397_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22603__B1 _15862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18851_ _13039_/B VGND VGND VPWR VPWR _18851_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24594__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17802_ _16678_/X _17798_/X _17801_/X VGND VGND VPWR VPWR _17802_/X sky130_fd_sc_hd__or3_4
XANTENNA__15636__A2 _15617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24523__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18782_ _18782_/A VGND VGND VPWR VPWR _18782_/Y sky130_fd_sc_hd__inv_2
X_15994_ _15991_/Y _15987_/X _15992_/X _15993_/X VGND VGND VPWR VPWR _15994_/X sky130_fd_sc_hd__a2bb2o_4
X_17733_ _17727_/A VGND VGND VPWR VPWR _17781_/A sky130_fd_sc_hd__buf_2
X_14945_ _15191_/A _22399_/A _15191_/A _22399_/A VGND VGND VPWR VPWR _14945_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17664_ _13406_/C _17663_/Y _17658_/X VGND VGND VPWR VPWR _17664_/X sky130_fd_sc_hd__o21a_4
X_14876_ _14876_/A _15034_/A _14876_/C _14876_/D VGND VGND VPWR VPWR _14877_/D sky130_fd_sc_hd__or4_4
X_19403_ _19401_/Y _19397_/X _19311_/X _19402_/X VGND VGND VPWR VPWR _23348_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16615_ _14818_/Y _16570_/A _16291_/X _16570_/A VGND VGND VPWR VPWR _24127_/D sky130_fd_sc_hd__a2bb2o_4
X_13827_ _13827_/A VGND VGND VPWR VPWR _13828_/D sky130_fd_sc_hd__buf_2
X_17595_ _16712_/Y _16700_/X _17595_/C _17607_/B VGND VGND VPWR VPWR _17595_/X sky130_fd_sc_hd__or4_4
XFILLER_16_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19334_ _19327_/Y VGND VGND VPWR VPWR _19334_/X sky130_fd_sc_hd__buf_2
XFILLER_1_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13758_ _13758_/A VGND VGND VPWR VPWR _13791_/A sky130_fd_sc_hd__inv_2
X_16546_ _16545_/X VGND VGND VPWR VPWR _16546_/X sky130_fd_sc_hd__buf_2
XFILLER_43_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12709_ _12609_/Y _12709_/B VGND VGND VPWR VPWR _12710_/D sky130_fd_sc_hd__or2_4
X_19265_ _19265_/A VGND VGND VPWR VPWR _19265_/Y sky130_fd_sc_hd__inv_2
X_13689_ _13677_/C VGND VGND VPWR VPWR _13689_/X sky130_fd_sc_hd__buf_2
X_16477_ _24188_/Q VGND VGND VPWR VPWR _16477_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21893__B2 _22218_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21856__A2_N _21838_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22782__B _22429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18216_ _18216_/A _18214_/Y _18167_/Y _18299_/B VGND VGND VPWR VPWR _18217_/C sky130_fd_sc_hd__or4_4
X_15428_ _21179_/A VGND VGND VPWR VPWR _15428_/X sky130_fd_sc_hd__buf_2
X_19196_ _19196_/A VGND VGND VPWR VPWR _19196_/X sky130_fd_sc_hd__buf_2
XANTENNA__19838__B2 _19831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15359_ _15358_/X VGND VGND VPWR VPWR _15359_/X sky130_fd_sc_hd__buf_2
X_18147_ _16075_/A _23864_/Q _16075_/Y _18205_/A VGND VGND VPWR VPWR _18154_/A sky130_fd_sc_hd__o22a_4
XFILLER_116_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17595__C _17595_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18078_ _18065_/C _18065_/B _18690_/B VGND VGND VPWR VPWR _18078_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16521__B1 _15369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17029_ _17028_/Y _17134_/A VGND VGND VPWR VPWR _17029_/X sky130_fd_sc_hd__or2_4
X_20040_ _20040_/A VGND VGND VPWR VPWR _21831_/B sky130_fd_sc_hd__inv_2
XFILLER_63_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22303__A _24478_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15088__B1 _14984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24264__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16301__A _16301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_70_0_HCLK clkbuf_8_71_0_HCLK/A VGND VGND VPWR VPWR _23789_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21991_ _22852_/A VGND VGND VPWR VPWR _21991_/X sky130_fd_sc_hd__buf_2
XFILLER_27_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23730_ _24349_/CLK _23730_/D HRESETn VGND VGND VPWR VPWR _23730_/Q sky130_fd_sc_hd__dfrtp_4
X_20942_ _21130_/A VGND VGND VPWR VPWR _22089_/A sky130_fd_sc_hd__buf_2
XFILLER_94_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16588__B1 _16259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20758__A _20861_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23661_ _23661_/CLK _20728_/X HRESETn VGND VGND VPWR VPWR _23661_/Q sky130_fd_sc_hd__dfrtp_4
X_20873_ _14264_/Y _20872_/X _14306_/A _15426_/X VGND VGND VPWR VPWR _20873_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17132__A _17132_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22612_ _22605_/X _22612_/B _22612_/C _22611_/X VGND VGND VPWR VPWR _22612_/X sky130_fd_sc_hd__or4_4
XPHY_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23592_ _23128_/CLK _23592_/D VGND VGND VPWR VPWR _13266_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14475__B _14437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16393__D _16393_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22543_ _12947_/A _20838_/X _17558_/B _22191_/X VGND VGND VPWR VPWR _22543_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25052__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22474_ _22474_/A _21978_/X VGND VGND VPWR VPWR _22474_/X sky130_fd_sc_hd__and2_4
X_24213_ _24213_/CLK _16417_/X HRESETn VGND VGND VPWR VPWR _24213_/Q sky130_fd_sc_hd__dfrtp_4
X_21425_ _16548_/Y _21425_/B VGND VGND VPWR VPWR _21425_/X sky130_fd_sc_hd__and2_4
XANTENNA__19059__A _18763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25193_ _23957_/CLK _25193_/D HRESETn VGND VGND VPWR VPWR _25193_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24144_ _24113_/CLK _16589_/X HRESETn VGND VGND VPWR VPWR _24144_/Q sky130_fd_sc_hd__dfrtp_4
X_21356_ _21339_/X _21355_/X _21175_/X VGND VGND VPWR VPWR _21356_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16512__B1 _16264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20307_ _18614_/X _20306_/Y _20315_/C VGND VGND VPWR VPWR _20307_/X sky130_fd_sc_hd__and3_4
X_24075_ _24079_/CLK _24075_/D HRESETn VGND VGND VPWR VPWR _24075_/Q sky130_fd_sc_hd__dfrtp_4
X_21287_ _22610_/A _21285_/X _21280_/X _21286_/X VGND VGND VPWR VPWR _21287_/X sky130_fd_sc_hd__o22a_4
XFILLER_1_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16741__A2_N _22979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23026_ _23026_/A _23026_/B VGND VGND VPWR VPWR _23026_/Y sky130_fd_sc_hd__nor2_4
X_20238_ _23694_/Q _20251_/B _20195_/X VGND VGND VPWR VPWR _20238_/X sky130_fd_sc_hd__a21o_4
XFILLER_118_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15618__A2 _15617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20169_ _20168_/B VGND VGND VPWR VPWR _20171_/B sky130_fd_sc_hd__buf_2
XFILLER_39_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12991_ _12863_/Y _12974_/B VGND VGND VPWR VPWR _12991_/Y sky130_fd_sc_hd__nand2_4
XFILLER_57_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13371__A1_N _13370_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24977_ _25141_/CLK _24977_/D HRESETn VGND VGND VPWR VPWR _24977_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11942_ _11941_/X VGND VGND VPWR VPWR _22616_/A sky130_fd_sc_hd__buf_2
X_14730_ _24706_/Q _24117_/Q _14868_/B _14729_/Y VGND VGND VPWR VPWR _14734_/C sky130_fd_sc_hd__o22a_4
XFILLER_57_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23928_ _23469_/CLK _23928_/D HRESETn VGND VGND VPWR VPWR _23928_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23987__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14661_ _24723_/Q _14612_/B _24723_/Q _14612_/B VGND VGND VPWR VPWR _14661_/X sky130_fd_sc_hd__a2bb2o_4
X_11873_ _11871_/B _11866_/X VGND VGND VPWR VPWR _11873_/X sky130_fd_sc_hd__and2_4
X_23859_ _23859_/CLK _18289_/Y HRESETn VGND VGND VPWR VPWR _23859_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23916__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13612_ _13612_/A VGND VGND VPWR VPWR _13613_/A sky130_fd_sc_hd__buf_2
X_16400_ _24219_/Q VGND VGND VPWR VPWR _16400_/Y sky130_fd_sc_hd__inv_2
X_14592_ _14553_/Y _14592_/B _18920_/A VGND VGND VPWR VPWR _14592_/X sky130_fd_sc_hd__and3_4
X_17380_ _17311_/Y _17371_/X VGND VGND VPWR VPWR _17380_/X sky130_fd_sc_hd__or2_4
XFILLER_60_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13543_ _23758_/Q _13543_/B VGND VGND VPWR VPWR _20551_/B sky130_fd_sc_hd__or2_4
X_16331_ _16330_/Y _16326_/X _16254_/X _16326_/X VGND VGND VPWR VPWR _16331_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16881__A _16858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16262_ _16262_/A VGND VGND VPWR VPWR _16262_/X sky130_fd_sc_hd__buf_2
X_19050_ _19048_/Y _19049_/X _18959_/X _19049_/X VGND VGND VPWR VPWR _19050_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21499__A _21235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13474_ _13474_/A _13474_/B _19946_/B _21257_/A VGND VGND VPWR VPWR _13480_/B sky130_fd_sc_hd__and4_4
XFILLER_72_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15213_ _15192_/A _15213_/B _15213_/C VGND VGND VPWR VPWR _24657_/D sky130_fd_sc_hd__and3_4
X_18001_ _17999_/X _17990_/X _18000_/X _23913_/Q _17974_/X VGND VGND VPWR VPWR _18001_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_9_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12425_ _12401_/X _12424_/X VGND VGND VPWR VPWR _12425_/X sky130_fd_sc_hd__or2_4
XANTENNA__12368__B2 _24480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15497__A HWDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16193_ _16193_/A VGND VGND VPWR VPWR _16193_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22824__B1 _24420_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15144_ _15144_/A _15144_/B _15143_/X VGND VGND VPWR VPWR _15144_/X sky130_fd_sc_hd__or3_4
XFILLER_103_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12356_ _12356_/A VGND VGND VPWR VPWR _12356_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24775__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15075_ _15057_/X _15075_/B _15075_/C VGND VGND VPWR VPWR _15075_/X sky130_fd_sc_hd__and3_4
X_19952_ _23148_/Q VGND VGND VPWR VPWR _19952_/Y sky130_fd_sc_hd__inv_2
X_12287_ _12122_/A _12287_/B VGND VGND VPWR VPWR _12288_/B sky130_fd_sc_hd__or2_4
XANTENNA__24704__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14026_ _14037_/B _14023_/X _14025_/Y VGND VGND VPWR VPWR _14026_/X sky130_fd_sc_hd__a21o_4
X_18903_ _17757_/B VGND VGND VPWR VPWR _18903_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19883_ _14493_/X _19883_/B _19883_/C VGND VGND VPWR VPWR _19883_/X sky130_fd_sc_hd__or3_4
XFILLER_45_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20063__B1 _15520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18834_ _22053_/B _18833_/X _15541_/X _18833_/X VGND VGND VPWR VPWR _23550_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11664__A2_N _23913_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16121__A _16121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_57_0_HCLK clkbuf_6_28_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_57_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18765_ _18758_/Y _18762_/X _18764_/X _18762_/X VGND VGND VPWR VPWR _23574_/D sky130_fd_sc_hd__a2bb2o_4
X_15977_ _22192_/A VGND VGND VPWR VPWR _15977_/Y sky130_fd_sc_hd__inv_2
X_17716_ _17726_/A VGND VGND VPWR VPWR _17716_/X sky130_fd_sc_hd__buf_2
XANTENNA__19432__A _19417_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14928_ _24668_/Q VGND VGND VPWR VPWR _15106_/A sky130_fd_sc_hd__inv_2
XFILLER_76_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18696_ _23596_/Q VGND VGND VPWR VPWR _18696_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21563__B1 _15395_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17647_ _21153_/A VGND VGND VPWR VPWR _21336_/A sky130_fd_sc_hd__buf_2
X_14859_ _14859_/A VGND VGND VPWR VPWR _14859_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23657__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13480__A _13480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17578_ _17494_/Y _17577_/X VGND VGND VPWR VPWR _17578_/X sky130_fd_sc_hd__or2_4
XFILLER_95_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19317_ _19316_/Y _19312_/X _19201_/X _19312_/X VGND VGND VPWR VPWR _19317_/X sky130_fd_sc_hd__a2bb2o_4
X_16529_ _24168_/Q VGND VGND VPWR VPWR _22282_/A sky130_fd_sc_hd__inv_2
XANTENNA__20669__A2 _13539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13630__D _22314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19248_ _23402_/Q VGND VGND VPWR VPWR _21484_/B sky130_fd_sc_hd__inv_2
XANTENNA__22815__B1 _24570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19179_ _23426_/Q VGND VGND VPWR VPWR _19179_/Y sky130_fd_sc_hd__inv_2
X_21210_ _21205_/A VGND VGND VPWR VPWR _21211_/A sky130_fd_sc_hd__buf_2
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22190_ _22163_/A _22189_/X VGND VGND VPWR VPWR _22190_/X sky130_fd_sc_hd__and2_4
XFILLER_121_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21141_ _21135_/X _21140_/X _18049_/X VGND VGND VPWR VPWR _21141_/X sky130_fd_sc_hd__o21a_4
XFILLER_105_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24445__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21072_ _21072_/A _21079_/B VGND VGND VPWR VPWR _21072_/X sky130_fd_sc_hd__or2_4
XFILLER_119_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20023_ _21605_/B _20020_/X _19721_/X _20020_/X VGND VGND VPWR VPWR _20023_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17127__A _24040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24900_ _24902_/CLK _13914_/X HRESETn VGND VGND VPWR VPWR _13810_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_112_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24831_ _24953_/CLK _24831_/D HRESETn VGND VGND VPWR VPWR MSO_S3 sky130_fd_sc_hd__dfrtp_4
XFILLER_80_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15481__B1 _11552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15870__A _24410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21591__B _21591_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24762_ _24968_/CLK _14406_/X HRESETn VGND VGND VPWR VPWR _24762_/Q sky130_fd_sc_hd__dfrtp_4
X_21974_ _22629_/A VGND VGND VPWR VPWR _21974_/X sky130_fd_sc_hd__buf_2
XANTENNA__20488__A _20465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23713_ _23716_/CLK _23713_/D HRESETn VGND VGND VPWR VPWR _20499_/B sky130_fd_sc_hd__dfrtp_4
X_20925_ _20925_/A VGND VGND VPWR VPWR _20925_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24693_ _24712_/CLK _24693_/D HRESETn VGND VGND VPWR VPWR _14694_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23644_ _23648_/CLK _23643_/Q HRESETn VGND VGND VPWR VPWR _23644_/Q sky130_fd_sc_hd__dfrtp_4
X_20856_ _20856_/A VGND VGND VPWR VPWR _21297_/A sky130_fd_sc_hd__inv_2
XFILLER_74_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23575_ _23568_/CLK _18757_/X VGND VGND VPWR VPWR _18756_/A sky130_fd_sc_hd__dfxtp_4
X_20787_ _24360_/Q _20787_/B VGND VGND VPWR VPWR _20787_/X sky130_fd_sc_hd__or2_4
XFILLER_126_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22526_ _21040_/X _22523_/Y _22260_/X _22525_/X VGND VGND VPWR VPWR _22526_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22457_ _22457_/A _22457_/B _22457_/C _22456_/X VGND VGND VPWR VPWR HRDATA[14] sky130_fd_sc_hd__or4_4
XFILLER_136_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ _25129_/Q _12214_/B VGND VGND VPWR VPWR _12210_/X sky130_fd_sc_hd__or2_4
XFILLER_108_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21408_ _24470_/Q _21408_/B VGND VGND VPWR VPWR _21408_/X sky130_fd_sc_hd__or2_4
X_13190_ _13222_/A _13184_/X _13190_/C VGND VGND VPWR VPWR _13191_/C sky130_fd_sc_hd__or3_4
XFILLER_109_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25176_ _23100_/CLK _25176_/D HRESETn VGND VGND VPWR VPWR _11826_/A sky130_fd_sc_hd__dfrtp_4
X_22388_ _16186_/A _22246_/B VGND VGND VPWR VPWR _22388_/X sky130_fd_sc_hd__or2_4
X_12141_ _25124_/Q VGND VGND VPWR VPWR _12171_/B sky130_fd_sc_hd__inv_2
XFILLER_123_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24127_ _24101_/CLK _24127_/D HRESETn VGND VGND VPWR VPWR _14818_/A sky130_fd_sc_hd__dfrtp_4
X_21339_ _21339_/A _21331_/X _21338_/X VGND VGND VPWR VPWR _21339_/X sky130_fd_sc_hd__or3_4
XANTENNA__24186__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23684__D _23684_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12072_ _12178_/C _24556_/Q _12178_/C _24556_/Q VGND VGND VPWR VPWR _12081_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24115__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24058_ _24612_/CLK _24058_/D HRESETn VGND VGND VPWR VPWR _24058_/Q sky130_fd_sc_hd__dfrtp_4
X_15900_ _15826_/A VGND VGND VPWR VPWR _15900_/X sky130_fd_sc_hd__buf_2
XFILLER_81_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23009_ _16621_/A _23008_/X _22839_/X _24576_/Q _21694_/X VGND VGND VPWR VPWR _23009_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17037__A _24039_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16880_ _16841_/D _16879_/X _16802_/Y VGND VGND VPWR VPWR _16880_/X sky130_fd_sc_hd__o21a_4
XFILLER_42_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15831_ _15830_/Y _15827_/X _11522_/X _15827_/X VGND VGND VPWR VPWR _24425_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21782__A _21224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16695__A2_N _20778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18550_ _18424_/D _18468_/C VGND VGND VPWR VPWR _18551_/B sky130_fd_sc_hd__or2_4
X_12974_ _12974_/A _12974_/B VGND VGND VPWR VPWR _12974_/X sky130_fd_sc_hd__or2_4
X_15762_ _12803_/Y _15757_/X _15761_/X _15757_/X VGND VGND VPWR VPWR _15762_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17501_ _17492_/X _17500_/X VGND VGND VPWR VPWR _17502_/D sky130_fd_sc_hd__or2_4
X_14713_ _24114_/Q VGND VGND VPWR VPWR _14713_/Y sky130_fd_sc_hd__inv_2
X_11925_ _21707_/A _11919_/X _11926_/A _11924_/X VGND VGND VPWR VPWR _11925_/X sky130_fd_sc_hd__a2bb2o_4
X_18481_ _18468_/B _18445_/X _18468_/A VGND VGND VPWR VPWR _18481_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15693_ _16581_/A VGND VGND VPWR VPWR _15693_/X sky130_fd_sc_hd__buf_2
XANTENNA__23750__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16567__A3 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17432_ _17321_/Y _17409_/B _17430_/B _17345_/X VGND VGND VPWR VPWR _17433_/A sky130_fd_sc_hd__a211o_4
XFILLER_2_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12038__B1 _11992_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11856_ _19617_/A VGND VGND VPWR VPWR _11856_/Y sky130_fd_sc_hd__inv_2
X_14644_ _14614_/C _14628_/X _14630_/A _14630_/B VGND VGND VPWR VPWR _14644_/X sky130_fd_sc_hd__o22a_4
XFILLER_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14575_ _17702_/A _14573_/X _14574_/Y VGND VGND VPWR VPWR _14575_/X sky130_fd_sc_hd__o21a_4
X_17363_ _17349_/B VGND VGND VPWR VPWR _17363_/Y sky130_fd_sc_hd__inv_2
X_11787_ _25184_/Q _11772_/B _11786_/Y VGND VGND VPWR VPWR _11787_/X sky130_fd_sc_hd__and3_4
X_19102_ _19099_/Y _19101_/X _19059_/X _19101_/X VGND VGND VPWR VPWR _19102_/X sky130_fd_sc_hd__a2bb2o_4
X_16314_ _16339_/A VGND VGND VPWR VPWR _16314_/X sky130_fd_sc_hd__buf_2
X_13526_ _13526_/A _13526_/B VGND VGND VPWR VPWR _13527_/B sky130_fd_sc_hd__nor2_4
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17294_ _11614_/Y _17239_/A _11628_/Y _17318_/A VGND VGND VPWR VPWR _17294_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24956__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22118__A _22198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19033_ _19799_/A _18072_/X _20134_/C VGND VGND VPWR VPWR _19034_/A sky130_fd_sc_hd__or3_4
X_13457_ _13474_/B VGND VGND VPWR VPWR _13458_/B sky130_fd_sc_hd__inv_2
X_16245_ _14956_/Y _16242_/X _15837_/X _16242_/X VGND VGND VPWR VPWR _24283_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12408_ _12344_/Y _12328_/Y _12408_/C _12408_/D VGND VGND VPWR VPWR _12505_/A sky130_fd_sc_hd__or4_4
XANTENNA__15020__A _15045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13388_ _20686_/B _13388_/B VGND VGND VPWR VPWR _13388_/X sky130_fd_sc_hd__and2_4
X_16176_ _24305_/Q VGND VGND VPWR VPWR _16176_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20861__A _15159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_20_0_HCLK clkbuf_4_10_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_41_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12339_ _24486_/Q VGND VGND VPWR VPWR _12339_/Y sky130_fd_sc_hd__inv_2
X_15127_ _14966_/Y _15125_/X _15126_/X _15119_/Y VGND VGND VPWR VPWR _15127_/X sky130_fd_sc_hd__a211o_4
XFILLER_99_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15955__A _22598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15058_ _15058_/A _14974_/X VGND VGND VPWR VPWR _15059_/B sky130_fd_sc_hd__or2_4
X_19935_ _21659_/B _19932_/X _19452_/A _19932_/X VGND VGND VPWR VPWR _23155_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22025__B2 _21868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14009_ _14009_/A VGND VGND VPWR VPWR _14009_/Y sky130_fd_sc_hd__inv_2
X_19866_ _23181_/Q VGND VGND VPWR VPWR _21956_/B sky130_fd_sc_hd__inv_2
XFILLER_110_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18817_ _16545_/X VGND VGND VPWR VPWR _18817_/X sky130_fd_sc_hd__buf_2
XFILLER_110_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19797_ _23207_/Q VGND VGND VPWR VPWR _19797_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23838__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22328__A2 _22230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18748_ _18747_/Y _18745_/X _18700_/X _18745_/X VGND VGND VPWR VPWR _18748_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22300__B _22246_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_144_0_HCLK clkbuf_7_72_0_HCLK/X VGND VGND VPWR VPWR _23128_/CLK sky130_fd_sc_hd__clkbuf_1
X_18679_ _18678_/X VGND VGND VPWR VPWR _18679_/X sky130_fd_sc_hd__buf_2
XFILLER_97_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20710_ _20710_/A _20710_/B _20710_/C VGND VGND VPWR VPWR _20710_/X sky130_fd_sc_hd__and3_4
X_21690_ _21689_/X VGND VGND VPWR VPWR _21705_/B sky130_fd_sc_hd__inv_2
X_20641_ _16508_/Y _20552_/X _20583_/X _20640_/Y VGND VGND VPWR VPWR _20642_/A sky130_fd_sc_hd__o22a_4
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23360_ _24998_/CLK _23360_/D VGND VGND VPWR VPWR _19365_/A sky130_fd_sc_hd__dfxtp_4
X_20572_ _16544_/Y _20553_/X _20562_/X _20571_/Y VGND VGND VPWR VPWR _20573_/A sky130_fd_sc_hd__o22a_4
XANTENNA__24697__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22311_ _22311_/A VGND VGND VPWR VPWR _22312_/B sky130_fd_sc_hd__buf_2
X_23291_ _23939_/CLK _23291_/D VGND VGND VPWR VPWR _23291_/Q sky130_fd_sc_hd__dfxtp_4
X_25030_ _24451_/CLK _12921_/X HRESETn VGND VGND VPWR VPWR _22826_/A sky130_fd_sc_hd__dfrtp_4
X_22242_ _21991_/X _22241_/X VGND VGND VPWR VPWR _22242_/X sky130_fd_sc_hd__and2_4
XFILLER_117_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21867__A _21867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22173_ _21069_/X VGND VGND VPWR VPWR _22173_/X sky130_fd_sc_hd__buf_2
X_21124_ _21124_/A _21590_/B VGND VGND VPWR VPWR _21124_/X sky130_fd_sc_hd__or2_4
XFILLER_117_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22016__B2 _22015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16788__A1_N _24396_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21055_ _21055_/A _21710_/B VGND VGND VPWR VPWR _21055_/X sky130_fd_sc_hd__or2_4
XFILLER_132_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22698__A _22698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20006_ _20005_/Y _20003_/X _19963_/X _20003_/X VGND VGND VPWR VPWR _23128_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_40_0_HCLK clkbuf_7_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_81_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24814_ _23774_/CLK _14233_/X HRESETn VGND VGND VPWR VPWR _14230_/A sky130_fd_sc_hd__dfstp_4
XFILLER_74_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21527__B1 _21242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21957_ _21378_/A _21957_/B VGND VGND VPWR VPWR _21957_/X sky130_fd_sc_hd__or2_4
XFILLER_76_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24745_ _25052_/CLK _14527_/X HRESETn VGND VGND VPWR VPWR _24745_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _13053_/C VGND VGND VPWR VPWR _11710_/X sky130_fd_sc_hd__buf_2
XANTENNA__11633__A _25192_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _17224_/Y _22497_/B _20903_/X _20907_/Y VGND VGND VPWR VPWR _20908_/X sky130_fd_sc_hd__a211o_4
X_12690_ _12571_/Y _12694_/B VGND VGND VPWR VPWR _12690_/Y sky130_fd_sc_hd__nand2_4
XPHY_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24676_ _24676_/CLK _15145_/Y HRESETn VGND VGND VPWR VPWR _24676_/Q sky130_fd_sc_hd__dfrtp_4
X_21888_ _21888_/A _22858_/A VGND VGND VPWR VPWR _21888_/X sky130_fd_sc_hd__and2_4
XPHY_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ HWDATA[0] VGND VGND VPWR VPWR _13644_/A sky130_fd_sc_hd__buf_2
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23627_ _23624_/CLK _20710_/B HRESETn VGND VGND VPWR VPWR _13923_/C sky130_fd_sc_hd__dfstp_4
X_20839_ _20838_/X VGND VGND VPWR VPWR _20839_/X sky130_fd_sc_hd__buf_2
XPHY_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _23651_/Q _14360_/B VGND VGND VPWR VPWR _14360_/X sky130_fd_sc_hd__and2_4
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ _25207_/Q VGND VGND VPWR VPWR _11572_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23041__B _20881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23558_ _24998_/CLK _18810_/X VGND VGND VPWR VPWR _13038_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_35_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ _13073_/A _13311_/B _13310_/X VGND VGND VPWR VPWR _13311_/X sky130_fd_sc_hd__or3_4
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22509_ _22879_/A _22502_/X _22504_/X _22507_/X _22508_/X VGND VGND VPWR VPWR _22509_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_7_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14291_ _14290_/Y _14288_/X _14232_/X _14288_/X VGND VGND VPWR VPWR _14291_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24367__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12464__A _12498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23489_ _23489_/CLK _19004_/X VGND VGND VPWR VPWR _19002_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22880__B _22806_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13242_ _13085_/A _19362_/A VGND VGND VPWR VPWR _13243_/C sky130_fd_sc_hd__or2_4
X_16030_ _24732_/Q _18759_/B _14587_/X VGND VGND VPWR VPWR _16030_/Y sky130_fd_sc_hd__o21ai_4
X_13173_ _13155_/X _13164_/X _13173_/C VGND VGND VPWR VPWR _13173_/X sky130_fd_sc_hd__and3_4
XFILLER_123_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15775__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25159_ _25159_/CLK _25159_/D HRESETn VGND VGND VPWR VPWR _11930_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_124_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12124_ _24546_/Q VGND VGND VPWR VPWR _12124_/Y sky130_fd_sc_hd__inv_2
X_17981_ _17999_/A VGND VGND VPWR VPWR _17982_/A sky130_fd_sc_hd__buf_2
XFILLER_111_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20018__B1 _19714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19720_ _23235_/Q VGND VGND VPWR VPWR _19720_/Y sky130_fd_sc_hd__inv_2
X_12055_ _25139_/Q _12053_/Y _12054_/X _12051_/A VGND VGND VPWR VPWR _12055_/X sky130_fd_sc_hd__a211o_4
X_16932_ _16936_/A _16932_/B _16931_/Y VGND VGND VPWR VPWR _24069_/D sky130_fd_sc_hd__and3_4
XFILLER_117_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17990__A _15430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19651_ _19651_/A VGND VGND VPWR VPWR _21832_/B sky130_fd_sc_hd__inv_2
X_16863_ _16863_/A _16769_/Y _16819_/Y _16874_/B VGND VGND VPWR VPWR _16866_/B sky130_fd_sc_hd__or4_4
XFILLER_77_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22401__A _22401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23931__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18602_ _18598_/X _18599_/X _18602_/C _18601_/X VGND VGND VPWR VPWR _18602_/X sky130_fd_sc_hd__or4_4
X_15814_ _15717_/X _15733_/X _15808_/X _15813_/X VGND VGND VPWR VPWR _15814_/X sky130_fd_sc_hd__a211o_4
XANTENNA__25155__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19582_ _21786_/B _19576_/X _19448_/X _19581_/X VGND VGND VPWR VPWR _19582_/X sky130_fd_sc_hd__a2bb2o_4
X_16794_ _15864_/Y _16784_/A _24416_/Q _16760_/Y VGND VGND VPWR VPWR _16796_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18533_ _18425_/A _18532_/X _18482_/A _18527_/Y VGND VGND VPWR VPWR _18534_/A sky130_fd_sc_hd__a211o_4
XFILLER_92_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15745_ _15744_/X VGND VGND VPWR VPWR _15746_/A sky130_fd_sc_hd__buf_2
X_12957_ _22474_/A _12957_/B VGND VGND VPWR VPWR _12959_/B sky130_fd_sc_hd__or2_4
XANTENNA__12639__A _12638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_217_0_HCLK clkbuf_7_108_0_HCLK/X VGND VGND VPWR VPWR _24213_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11908_ _11904_/Y _20691_/A _11904_/Y _20691_/A VGND VGND VPWR VPWR _11916_/B sky130_fd_sc_hd__a2bb2o_4
X_18464_ _18475_/A VGND VGND VPWR VPWR _18482_/A sky130_fd_sc_hd__buf_2
X_15676_ _12384_/Y _15669_/X _11558_/X _15669_/X VGND VGND VPWR VPWR _15676_/X sky130_fd_sc_hd__a2bb2o_4
X_12888_ _12890_/B VGND VGND VPWR VPWR _12888_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17415_ _17415_/A _17421_/B VGND VGND VPWR VPWR _17419_/B sky130_fd_sc_hd__or2_4
XFILLER_18_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14627_ _14612_/C _14627_/B _24725_/Q VGND VGND VPWR VPWR _14627_/X sky130_fd_sc_hd__or3_4
X_11839_ _19600_/A VGND VGND VPWR VPWR _11839_/X sky130_fd_sc_hd__buf_2
X_18395_ _23841_/Q VGND VGND VPWR VPWR _18452_/C sky130_fd_sc_hd__inv_2
X_17346_ _17340_/A _17339_/X _17345_/X _17342_/B VGND VGND VPWR VPWR _17347_/A sky130_fd_sc_hd__a211o_4
XFILLER_105_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18698__B1 _17205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14558_ _17674_/A _17877_/A VGND VGND VPWR VPWR _14558_/X sky130_fd_sc_hd__and2_4
XANTENNA__24790__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24811__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13509_ _13509_/A _13509_/B _13509_/C VGND VGND VPWR VPWR _13509_/X sky130_fd_sc_hd__or3_4
XFILLER_53_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17277_ _17277_/A _17274_/X _17277_/C _17277_/D VGND VGND VPWR VPWR _17277_/X sky130_fd_sc_hd__or4_4
X_14489_ _24741_/Q _14460_/X VGND VGND VPWR VPWR _14489_/X sky130_fd_sc_hd__and2_4
X_19016_ _21946_/B _19013_/X _15545_/X _19013_/X VGND VGND VPWR VPWR _23485_/D sky130_fd_sc_hd__a2bb2o_4
X_16228_ _16228_/A VGND VGND VPWR VPWR _16228_/X sky130_fd_sc_hd__buf_2
XANTENNA__24037__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14723__A2 _14722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15685__A _15664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16159_ _16157_/Y _16152_/X _15761_/X _16158_/X VGND VGND VPWR VPWR _24313_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18061__A _17446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16476__A2 _15415_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19918_ _19918_/A VGND VGND VPWR VPWR _19918_/X sky130_fd_sc_hd__buf_2
XFILLER_114_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19849_ _23187_/Q VGND VGND VPWR VPWR _21669_/B sky130_fd_sc_hd__inv_2
XANTENNA__22311__A _22311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23672__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_27_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22860_ _24281_/Q _22859_/X _22338_/A VGND VGND VPWR VPWR _22860_/X sky130_fd_sc_hd__o21a_4
X_21811_ _20972_/A _19538_/Y VGND VGND VPWR VPWR _21811_/X sky130_fd_sc_hd__or2_4
XFILLER_3_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17124__B _17124_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22791_ _22791_/A VGND VGND VPWR VPWR _22800_/C sky130_fd_sc_hd__inv_2
XFILLER_52_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22721__A2 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24530_ _25005_/CLK _15592_/X HRESETn VGND VGND VPWR VPWR _24530_/Q sky130_fd_sc_hd__dfrtp_4
X_21742_ _14272_/Y _21408_/B _24789_/Q _21400_/A VGND VGND VPWR VPWR _21742_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15739__A1 _15411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20732__A1 _23660_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24878__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24461_ _24944_/CLK _15742_/X HRESETn VGND VGND VPWR VPWR _24461_/Q sky130_fd_sc_hd__dfrtp_4
X_21673_ _21657_/A _21673_/B VGND VGND VPWR VPWR _21675_/B sky130_fd_sc_hd__or2_4
XFILLER_71_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23412_ _25194_/CLK _19219_/X VGND VGND VPWR VPWR _23412_/Q sky130_fd_sc_hd__dfxtp_4
X_20624_ _20651_/A VGND VGND VPWR VPWR _20624_/X sky130_fd_sc_hd__buf_2
XFILLER_71_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24392_ _24071_/CLK _15917_/X HRESETn VGND VGND VPWR VPWR _24392_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14483__B _14482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17497__D _17497_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23343_ _23343_/CLK _23343_/D VGND VGND VPWR VPWR _13313_/B sky130_fd_sc_hd__dfxtp_4
X_20555_ _20555_/A VGND VGND VPWR VPWR _20647_/A sky130_fd_sc_hd__buf_2
XANTENNA__24460__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15911__A1 _11535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23274_ _23258_/CLK _19611_/X VGND VGND VPWR VPWR _23274_/Q sky130_fd_sc_hd__dfxtp_4
X_20486_ _20517_/A VGND VGND VPWR VPWR _20495_/B sky130_fd_sc_hd__inv_2
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25013_ _24435_/CLK _12988_/X HRESETn VGND VGND VPWR VPWR _22160_/A sky130_fd_sc_hd__dfrtp_4
X_22225_ _22225_/A VGND VGND VPWR VPWR _22225_/X sky130_fd_sc_hd__buf_2
XANTENNA__22788__A2 _22170_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21996__B1 _11614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22156_ _16454_/Y _15572_/A _21715_/X _22155_/X VGND VGND VPWR VPWR _22157_/A sky130_fd_sc_hd__a211o_4
XFILLER_65_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_109_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_219_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21107_ _21106_/X VGND VGND VPWR VPWR _21107_/X sky130_fd_sc_hd__buf_2
XFILLER_133_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11628__A _25193_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22087_ _22087_/A _22087_/B VGND VGND VPWR VPWR _22089_/B sky130_fd_sc_hd__or2_4
XFILLER_102_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21038_ _21029_/X _21038_/B VGND VGND VPWR VPWR _21038_/X sky130_fd_sc_hd__and2_4
XANTENNA__15690__A3 _16093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22960__A2 _21576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13860_ _13869_/A _13830_/C VGND VGND VPWR VPWR _13872_/A sky130_fd_sc_hd__or2_4
X_12811_ _22651_/A _22633_/A _12809_/Y _12810_/Y VGND VGND VPWR VPWR _12811_/X sky130_fd_sc_hd__o22a_4
X_13791_ _13791_/A _14071_/D _13777_/X _13790_/X VGND VGND VPWR VPWR _13792_/C sky130_fd_sc_hd__or4_4
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22989_ _16310_/A _15919_/X _22858_/X _22988_/X VGND VGND VPWR VPWR _22990_/C sky130_fd_sc_hd__a211o_4
X_15530_ _15421_/X _15319_/Y _15432_/X _20413_/A _15529_/X VGND VGND VPWR VPWR _15530_/X
+ sky130_fd_sc_hd__a32o_4
X_12742_ _12581_/Y _12742_/B VGND VGND VPWR VPWR _12742_/X sky130_fd_sc_hd__or2_4
X_24728_ _24728_/CLK _24728_/D HRESETn VGND VGND VPWR VPWR _14614_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_31_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_190_0_HCLK clkbuf_7_95_0_HCLK/X VGND VGND VPWR VPWR _25084_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__23052__A _23036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12673_ _12637_/X _12673_/B _12673_/C VGND VGND VPWR VPWR _25066_/D sky130_fd_sc_hd__and3_4
X_15461_ _15460_/X VGND VGND VPWR VPWR _15461_/X sky130_fd_sc_hd__buf_2
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24548__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24659_ _24662_/CLK _15209_/X HRESETn VGND VGND VPWR VPWR _24659_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _20401_/A _17198_/X _17199_/X _17198_/X VGND VGND VPWR VPWR _24019_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_47_0_HCLK clkbuf_8_47_0_HCLK/A VGND VGND VPWR VPWR _23133_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ HWDATA[4] VGND VGND VPWR VPWR _11625_/A sky130_fd_sc_hd__buf_2
X_14412_ _14390_/D VGND VGND VPWR VPWR _14412_/X sky130_fd_sc_hd__buf_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17050__A _24058_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ _16116_/Y _23849_/Q _16054_/A _18179_/Y VGND VGND VPWR VPWR _18180_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ _24589_/Q VGND VGND VPWR VPWR _21728_/A sky130_fd_sc_hd__inv_2
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17131_ _17131_/A VGND VGND VPWR VPWR _17131_/Y sky130_fd_sc_hd__inv_2
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11555_ HWDATA[23] VGND VGND VPWR VPWR _11555_/X sky130_fd_sc_hd__buf_2
X_14343_ _14335_/X _14342_/X _24786_/Q _14320_/Y VGND VGND VPWR VPWR _14343_/X sky130_fd_sc_hd__o22a_4
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14274_ _14272_/Y _14268_/X _14236_/X _14273_/X VGND VGND VPWR VPWR _24797_/D sky130_fd_sc_hd__a2bb2o_4
X_17062_ _24056_/Q _17062_/B VGND VGND VPWR VPWR _17064_/B sky130_fd_sc_hd__or2_4
XANTENNA__24130__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13225_ _13057_/X _13224_/X _24999_/Q _13116_/X VGND VGND VPWR VPWR _24999_/D sky130_fd_sc_hd__o22a_4
X_16013_ _16012_/X VGND VGND VPWR VPWR _16014_/C sky130_fd_sc_hd__inv_2
XANTENNA__21300__A _21300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12922__A _12922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13156_ _13297_/A _13156_/B VGND VGND VPWR VPWR _13156_/X sky130_fd_sc_hd__or2_4
XANTENNA__21451__A2 _15653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12107_ _25131_/Q VGND VGND VPWR VPWR _12170_/A sky130_fd_sc_hd__inv_2
X_13087_ _13207_/A _13087_/B _13087_/C VGND VGND VPWR VPWR _13088_/C sky130_fd_sc_hd__or3_4
X_17964_ _17861_/A _18917_/A VGND VGND VPWR VPWR _17965_/C sky130_fd_sc_hd__or2_4
XANTENNA__21954__B _19783_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16618__A1_N _16616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19703_ _23240_/Q VGND VGND VPWR VPWR _19703_/Y sky130_fd_sc_hd__inv_2
X_12038_ _11992_/Y _20698_/A _11992_/Y _20698_/A VGND VGND VPWR VPWR _12045_/B sky130_fd_sc_hd__a2bb2o_4
X_16915_ _16829_/A _16915_/B VGND VGND VPWR VPWR _16917_/B sky130_fd_sc_hd__or2_4
XANTENNA__22400__A1 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22400__B2 _22228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17895_ _17895_/A _19091_/A VGND VGND VPWR VPWR _17895_/X sky130_fd_sc_hd__or2_4
XFILLER_38_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19634_ _21469_/B _19629_/X _19610_/X _19629_/X VGND VGND VPWR VPWR _23266_/D sky130_fd_sc_hd__a2bb2o_4
X_16846_ _16846_/A _16844_/Y VGND VGND VPWR VPWR _16846_/Y sky130_fd_sc_hd__nand2_4
XFILLER_93_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16091__B1 _11585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21970__A _21256_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19565_ _21477_/B _19560_/X _11853_/X _19560_/X VGND VGND VPWR VPWR _23290_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16777_ _24404_/Q _16776_/A _15884_/Y _16927_/A VGND VGND VPWR VPWR _16782_/B sky130_fd_sc_hd__o22a_4
X_13989_ _24884_/Q _13926_/B _24884_/Q _13926_/B VGND VGND VPWR VPWR _13989_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18516_ _18518_/B VGND VGND VPWR VPWR _18517_/B sky130_fd_sc_hd__inv_2
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15728_ _15728_/A VGND VGND VPWR VPWR _15729_/A sky130_fd_sc_hd__inv_2
X_19496_ _23315_/Q VGND VGND VPWR VPWR _21654_/B sky130_fd_sc_hd__inv_2
XANTENNA__20714__A1 _23622_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24971__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18447_ _18440_/B _18446_/X VGND VGND VPWR VPWR _18447_/X sky130_fd_sc_hd__or2_4
X_15659_ _16305_/A _15659_/B VGND VGND VPWR VPWR _15664_/A sky130_fd_sc_hd__or2_4
XANTENNA__24289__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24900__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21074__A1_N _14004_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18378_ _18347_/X _18378_/B _18367_/X _18377_/X VGND VGND VPWR VPWR _18378_/X sky130_fd_sc_hd__or4_4
XANTENNA__24218__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17329_ _17329_/A _17260_/Y _17340_/A _17328_/X VGND VGND VPWR VPWR _17329_/X sky130_fd_sc_hd__or4_4
XFILLER_119_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20340_ _20189_/A _20192_/X _13916_/X VGND VGND VPWR VPWR _23649_/D sky130_fd_sc_hd__o21a_4
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20271_ _20271_/A _13916_/X _13842_/X VGND VGND VPWR VPWR _23620_/D sky130_fd_sc_hd__and3_4
XFILLER_115_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19096__B1 _19095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11526__A1_N _11524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22010_ _21886_/X _22009_/X VGND VGND VPWR VPWR _22010_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__23853__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25077__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25006__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23961_ _23949_/CLK _17560_/X HRESETn VGND VGND VPWR VPWR _23961_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22041__A _21582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13663__A _13663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22942__A2 _22940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22912_ _22971_/A _22911_/X VGND VGND VPWR VPWR _22912_/X sky130_fd_sc_hd__and2_4
X_23892_ _23990_/CLK _18084_/X HRESETn VGND VGND VPWR VPWR _11733_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22843_ _13358_/X VGND VGND VPWR VPWR _23026_/B sky130_fd_sc_hd__buf_2
XFILLER_37_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22695__B _22435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19350__A _19349_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22774_ _22201_/A _22759_/X _22762_/X _22768_/X _22773_/X VGND VGND VPWR VPWR _22775_/D
+ sky130_fd_sc_hd__o41a_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_200_0_HCLK clkbuf_8_201_0_HCLK/A VGND VGND VPWR VPWR _24031_/CLK sky130_fd_sc_hd__clkbuf_1
X_21725_ _11999_/Y _11954_/X _24098_/Q _21570_/A VGND VGND VPWR VPWR _21725_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24513_ _24432_/CLK _24513_/D HRESETn VGND VGND VPWR VPWR _24513_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24641__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_6_0_HCLK clkbuf_8_7_0_HCLK/A VGND VGND VPWR VPWR _23258_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21656_ _21237_/A _21654_/X _21655_/X VGND VGND VPWR VPWR _21656_/X sky130_fd_sc_hd__and3_4
X_24444_ _24445_/CLK _24444_/D HRESETn VGND VGND VPWR VPWR _22463_/A sky130_fd_sc_hd__dfrtp_4
X_20607_ _20605_/Y _20599_/Y _20606_/X VGND VGND VPWR VPWR _20607_/X sky130_fd_sc_hd__o21a_4
X_24375_ _24385_/CLK _15964_/X HRESETn VGND VGND VPWR VPWR _22458_/A sky130_fd_sc_hd__dfrtp_4
X_21587_ _21300_/A _12061_/B _21587_/C VGND VGND VPWR VPWR _21587_/X sky130_fd_sc_hd__and3_4
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23326_ _24748_/CLK _19469_/X VGND VGND VPWR VPWR _23326_/Q sky130_fd_sc_hd__dfxtp_4
X_20538_ _20542_/B _13514_/X VGND VGND VPWR VPWR _20538_/Y sky130_fd_sc_hd__nor2_4
XFILLER_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21120__A SSn_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19087__B1 _18953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23257_ _23385_/CLK _23257_/D VGND VGND VPWR VPWR _23257_/Q sky130_fd_sc_hd__dfxtp_4
X_20469_ _20468_/A _20469_/B VGND VGND VPWR VPWR _20469_/X sky130_fd_sc_hd__or2_4
X_13010_ _13009_/Y _12921_/A _24461_/Q VGND VGND VPWR VPWR _25004_/D sky130_fd_sc_hd__a21oi_4
XFILLER_134_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22208_ _11913_/Y _21707_/B _16450_/A _22931_/A VGND VGND VPWR VPWR _22208_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22630__A1 _22116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21433__A2 _21292_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22630__B2 _22118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23188_ _23179_/CLK _23188_/D VGND VGND VPWR VPWR _23188_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20641__B1 _20583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22139_ _16534_/Y _22011_/X _15383_/Y _20927_/X VGND VGND VPWR VPWR _22139_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15663__A3 _15468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14961_ _24670_/Q VGND VGND VPWR VPWR _15161_/A sky130_fd_sc_hd__inv_2
XFILLER_59_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16700_ _16700_/A VGND VGND VPWR VPWR _16700_/X sky130_fd_sc_hd__buf_2
X_13912_ _13808_/X _13908_/X _13905_/X _13806_/X _13911_/X VGND VGND VPWR VPWR _13912_/X
+ sky130_fd_sc_hd__a32o_4
X_17680_ _17673_/X _17679_/X _16678_/X VGND VGND VPWR VPWR _17680_/X sky130_fd_sc_hd__o21a_4
X_14892_ _15138_/A _24280_/Q _14890_/Y _24280_/Q VGND VGND VPWR VPWR _14893_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22886__A _22885_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16631_ _14777_/Y _16629_/X _11536_/X _16629_/X VGND VGND VPWR VPWR _24121_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_10_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_13843_ _24899_/Q _24898_/Q VGND VGND VPWR VPWR _13843_/Y sky130_fd_sc_hd__nand2_4
XFILLER_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24729__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19350_ _19349_/Y VGND VGND VPWR VPWR _19350_/X sky130_fd_sc_hd__buf_2
X_16562_ _21590_/B VGND VGND VPWR VPWR _20863_/A sky130_fd_sc_hd__buf_2
XANTENNA__22697__A1 _22011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13774_ _13780_/B _13774_/B VGND VGND VPWR VPWR _13777_/C sky130_fd_sc_hd__nor2_4
X_18301_ _18214_/Y _18301_/B VGND VGND VPWR VPWR _18321_/A sky130_fd_sc_hd__or2_4
X_15513_ HWDATA[8] VGND VGND VPWR VPWR _15513_/X sky130_fd_sc_hd__buf_2
X_12725_ _12725_/A VGND VGND VPWR VPWR _12725_/Y sky130_fd_sc_hd__inv_2
X_19281_ _23390_/Q VGND VGND VPWR VPWR _22103_/B sky130_fd_sc_hd__inv_2
X_16493_ _16493_/A VGND VGND VPWR VPWR _16493_/X sky130_fd_sc_hd__buf_2
XANTENNA__24382__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18232_ _18179_/Y _18231_/X VGND VGND VPWR VPWR _18232_/X sky130_fd_sc_hd__or2_4
XFILLER_30_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15444_ _15443_/X VGND VGND VPWR VPWR _15449_/B sky130_fd_sc_hd__inv_2
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24311__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12656_ _12547_/Y _12679_/C _12655_/X VGND VGND VPWR VPWR _12663_/A sky130_fd_sc_hd__or3_4
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11607_ HWDATA[8] VGND VGND VPWR VPWR _11607_/X sky130_fd_sc_hd__buf_2
X_18163_ _18163_/A _18158_/X _18160_/X _18163_/D VGND VGND VPWR VPWR _18163_/X sky130_fd_sc_hd__or4_4
XFILLER_129_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12587_ _25055_/Q VGND VGND VPWR VPWR _12587_/Y sky130_fd_sc_hd__inv_2
X_15375_ _22344_/A _15366_/X _11594_/X _15374_/X VGND VGND VPWR VPWR _15375_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21121__A1 SSn_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17114_ _17042_/D _17096_/B _17083_/X _17112_/B VGND VGND VPWR VPWR _17115_/A sky130_fd_sc_hd__a211o_4
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14326_ _24780_/Q VGND VGND VPWR VPWR _14326_/Y sky130_fd_sc_hd__inv_2
X_11538_ _11533_/X _11535_/X _11536_/X _25218_/Q _11537_/X VGND VGND VPWR VPWR _11538_/X
+ sky130_fd_sc_hd__a32o_4
X_18094_ _18091_/Y _11767_/X _18093_/Y VGND VGND VPWR VPWR _18104_/B sky130_fd_sc_hd__o21ai_4
XFILLER_128_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17045_ _17077_/A _17076_/A _17045_/C _17044_/X VGND VGND VPWR VPWR _17045_/X sky130_fd_sc_hd__or4_4
XFILLER_99_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14257_ _14257_/A VGND VGND VPWR VPWR _14257_/Y sky130_fd_sc_hd__inv_2
X_13208_ _13155_/X _13200_/X _13208_/C VGND VGND VPWR VPWR _13208_/X sky130_fd_sc_hd__and3_4
XANTENNA__22621__A1 _16075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14188_ _24826_/Q _14169_/B _24825_/Q _14165_/B VGND VGND VPWR VPWR _14188_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21975__A3 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25170__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13139_ _13299_/A VGND VGND VPWR VPWR _13278_/A sky130_fd_sc_hd__buf_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18996_ _18990_/Y VGND VGND VPWR VPWR _18996_/X sky130_fd_sc_hd__buf_2
XFILLER_135_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17947_ _17947_/A _17943_/X _17947_/C VGND VGND VPWR VPWR _17947_/X sky130_fd_sc_hd__or3_4
XFILLER_100_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17878_ _17878_/A _19136_/A VGND VGND VPWR VPWR _17879_/C sky130_fd_sc_hd__or2_4
X_16829_ _16829_/A VGND VGND VPWR VPWR _16916_/A sky130_fd_sc_hd__inv_2
X_19617_ _19617_/A VGND VGND VPWR VPWR _19617_/X sky130_fd_sc_hd__buf_2
XFILLER_81_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19170__A _18763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19548_ _23296_/Q VGND VGND VPWR VPWR _19548_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22152__A3 _22150_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19479_ _23321_/Q VGND VGND VPWR VPWR _19479_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12827__A _21851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21510_ _21394_/A _21508_/X _21509_/X VGND VGND VPWR VPWR _21510_/X sky130_fd_sc_hd__and3_4
X_22490_ _22407_/X _22490_/B VGND VGND VPWR VPWR _22490_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24052__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_30_0_HCLK clkbuf_8_31_0_HCLK/A VGND VGND VPWR VPWR _23109_/CLK sky130_fd_sc_hd__clkbuf_1
X_21441_ _13326_/A _21439_/X _11954_/A _21440_/X VGND VGND VPWR VPWR _21441_/X sky130_fd_sc_hd__o22a_4
XFILLER_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21112__A1 _20926_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18514__A _18468_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_93_0_HCLK clkbuf_8_93_0_HCLK/A VGND VGND VPWR VPWR _23664_/CLK sky130_fd_sc_hd__clkbuf_1
X_24160_ _24161_/CLK _24160_/D HRESETn VGND VGND VPWR VPWR _24160_/Q sky130_fd_sc_hd__dfrtp_4
X_21372_ _21372_/A _21372_/B _21372_/C VGND VGND VPWR VPWR _21372_/X sky130_fd_sc_hd__and3_4
XFILLER_119_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22860__A1 _24281_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15878__B1 _11594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23111_ _23112_/CLK _23111_/D VGND VGND VPWR VPWR _23111_/Q sky130_fd_sc_hd__dfxtp_4
X_20323_ _18619_/B VGND VGND VPWR VPWR _20323_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13658__A _15788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19069__B1 _18932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24091_ _24071_/CLK _16750_/X HRESETn VGND VGND VPWR VPWR _20737_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_134_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23042_ _25156_/Q _23042_/B VGND VGND VPWR VPWR _23042_/X sky130_fd_sc_hd__and2_4
X_20254_ _20254_/A _23773_/Q _20244_/A _20254_/D VGND VGND VPWR VPWR _20254_/X sky130_fd_sc_hd__or4_4
XFILLER_116_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16969__A _24054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20185_ _20185_/A _20184_/Y VGND VGND VPWR VPWR _20185_/Y sky130_fd_sc_hd__nor2_4
XFILLER_89_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21594__B _13333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24993_ _24841_/CLK _13342_/X HRESETn VGND VGND VPWR VPWR _13341_/A sky130_fd_sc_hd__dfrtp_4
X_23944_ _23972_/CLK _23944_/D HRESETn VGND VGND VPWR VPWR _23944_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12864__B1 _12858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24893__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16055__B1 _15837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24822__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23875_ _23767_/CLK _18230_/Y HRESETn VGND VGND VPWR VPWR _23875_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15802__B1 _15801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22826_ _22826_/A _22651_/B VGND VGND VPWR VPWR _22826_/X sky130_fd_sc_hd__and2_4
XFILLER_129_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12092__B2 _24545_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22757_ _24490_/Q _22757_/B VGND VGND VPWR VPWR _22757_/X sky130_fd_sc_hd__or2_4
XANTENNA__11641__A HWDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12510_ _12408_/C _12505_/B VGND VGND VPWR VPWR _12511_/D sky130_fd_sc_hd__or2_4
X_13490_ _13488_/X _13490_/B VGND VGND VPWR VPWR _13490_/X sky130_fd_sc_hd__or2_4
X_21708_ _18117_/Y _11954_/X _17134_/A _20747_/X VGND VGND VPWR VPWR _21708_/X sky130_fd_sc_hd__o22a_4
XFILLER_12_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14908__A2 _24274_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22688_ _24114_/Q _22574_/B VGND VGND VPWR VPWR _22688_/X sky130_fd_sc_hd__or2_4
X_12441_ _12434_/A _12439_/X _12440_/X VGND VGND VPWR VPWR _25097_/D sky130_fd_sc_hd__and3_4
X_21639_ _20062_/Y _21638_/X _20122_/Y _21795_/B VGND VGND VPWR VPWR _21639_/X sky130_fd_sc_hd__o22a_4
XFILLER_12_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24427_ _23442_/CLK _15817_/X HRESETn VGND VGND VPWR VPWR _15713_/A sky130_fd_sc_hd__dfrtp_4
X_12372_ _12412_/B _22565_/A _12469_/A _12319_/Y VGND VGND VPWR VPWR _12376_/C sky130_fd_sc_hd__a2bb2o_4
X_15160_ _15107_/C _15159_/X VGND VGND VPWR VPWR _15161_/B sky130_fd_sc_hd__or2_4
XFILLER_138_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24358_ _25183_/CLK _24358_/D HRESETn VGND VGND VPWR VPWR _16014_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23775__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_1_0_HCLK clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__15869__B1 _11576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14111_ _14107_/Y _14108_/Y _14111_/C _14110_/X VGND VGND VPWR VPWR _14111_/X sky130_fd_sc_hd__or4_4
XFILLER_138_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15091_ _14867_/A _15087_/X _15090_/Y VGND VGND VPWR VPWR _15091_/X sky130_fd_sc_hd__and3_4
X_23309_ _23282_/CLK _23309_/D VGND VGND VPWR VPWR _23309_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24289_ _24289_/CLK _24289_/D HRESETn VGND VGND VPWR VPWR _24289_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23704__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14042_ _20719_/A _14037_/X _13645_/X _14027_/X VGND VGND VPWR VPWR _14042_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18850_ _18849_/Y _18845_/X _18662_/X _18832_/Y VGND VGND VPWR VPWR _23543_/D sky130_fd_sc_hd__a2bb2o_4
X_17801_ _14569_/A _17799_/X _17800_/X VGND VGND VPWR VPWR _17801_/X sky130_fd_sc_hd__and3_4
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15636__A3 _15635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18781_ _18780_/Y _18776_/X _18712_/X _18776_/A VGND VGND VPWR VPWR _23567_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15993_ _15921_/X VGND VGND VPWR VPWR _15993_/X sky130_fd_sc_hd__buf_2
XANTENNA__22367__B1 _24514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17732_ _17732_/A VGND VGND VPWR VPWR _17783_/A sky130_fd_sc_hd__buf_2
XFILLER_48_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14944_ _15190_/A VGND VGND VPWR VPWR _15191_/A sky130_fd_sc_hd__inv_2
XFILLER_76_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12855__B1 _12854_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17663_ _17663_/A VGND VGND VPWR VPWR _17663_/Y sky130_fd_sc_hd__inv_2
X_14875_ _14770_/Y _14759_/Y _14874_/Y _15022_/A VGND VGND VPWR VPWR _14875_/X sky130_fd_sc_hd__or4_4
XANTENNA__22119__B1 _25197_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24563__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19402_ _19396_/Y VGND VGND VPWR VPWR _19402_/X sky130_fd_sc_hd__buf_2
XFILLER_29_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16614_ _15657_/X _16597_/X _15706_/X _24128_/Q _16590_/X VGND VGND VPWR VPWR _24128_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_62_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13826_ _13818_/A VGND VGND VPWR VPWR _13828_/C sky130_fd_sc_hd__buf_2
X_17594_ _16685_/Y _17594_/B VGND VGND VPWR VPWR _17607_/B sky130_fd_sc_hd__or2_4
XFILLER_1_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19333_ _19333_/A VGND VGND VPWR VPWR _19333_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19535__B2 _19534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16545_ HWDATA[4] VGND VGND VPWR VPWR _16545_/X sky130_fd_sc_hd__buf_2
XFILLER_90_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13757_ _13757_/A _13757_/B _13769_/C _13782_/B VGND VGND VPWR VPWR _13758_/A sky130_fd_sc_hd__or4_4
X_12708_ _12644_/D _12700_/B VGND VGND VPWR VPWR _12709_/B sky130_fd_sc_hd__or2_4
X_19264_ _19263_/Y _19261_/X _19149_/X _19261_/X VGND VGND VPWR VPWR _23397_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16476_ _15619_/X _15415_/Y _15743_/X _24189_/Q _16475_/X VGND VGND VPWR VPWR _24189_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21893__A2 _21300_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13688_ _20201_/B VGND VGND VPWR VPWR _13688_/Y sky130_fd_sc_hd__inv_2
X_18215_ _23845_/Q VGND VGND VPWR VPWR _18299_/B sky130_fd_sc_hd__inv_2
X_15427_ _15426_/X VGND VGND VPWR VPWR _21179_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_17_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_12639_ _12638_/Y VGND VGND VPWR VPWR _12727_/A sky130_fd_sc_hd__buf_2
X_19195_ _23420_/Q VGND VGND VPWR VPWR _19195_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18146_ _23864_/Q VGND VGND VPWR VPWR _18205_/A sky130_fd_sc_hd__inv_2
X_15358_ _15401_/A VGND VGND VPWR VPWR _15358_/X sky130_fd_sc_hd__buf_2
XFILLER_15_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14309_ _20164_/B VGND VGND VPWR VPWR _14309_/X sky130_fd_sc_hd__buf_2
X_18077_ _19303_/A _18690_/B _19303_/A _18690_/B VGND VGND VPWR VPWR _23895_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15289_ _15288_/Y _15285_/X _14304_/X _15285_/X VGND VGND VPWR VPWR _24626_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17028_ _24038_/Q VGND VGND VPWR VPWR _17028_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15693__A _16581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19471__B1 _19421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16285__B1 _15894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22303__B _22999_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18979_ _13197_/B VGND VGND VPWR VPWR _18979_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16301__B _22230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11726__A _11725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21990_ _21990_/A VGND VGND VPWR VPWR _22852_/A sky130_fd_sc_hd__buf_2
XANTENNA__20908__A1 _17224_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12846__B1 _22258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20941_ _23939_/Q VGND VGND VPWR VPWR _21130_/A sky130_fd_sc_hd__buf_2
XFILLER_96_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20872_ _11500_/X VGND VGND VPWR VPWR _20872_/X sky130_fd_sc_hd__buf_2
XFILLER_82_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24233__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23660_ _24643_/CLK _23660_/D HRESETn VGND VGND VPWR VPWR _23660_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22611_ _20498_/Y _22610_/X _20635_/B _22531_/X VGND VGND VPWR VPWR _22611_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23591_ _23596_/CLK _18713_/X VGND VGND VPWR VPWR _23591_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12074__B2 _24576_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22542_ _22943_/A _22541_/X VGND VGND VPWR VPWR _22542_/Y sky130_fd_sc_hd__nor2_4
X_22473_ _22473_/A _22256_/B VGND VGND VPWR VPWR _22473_/X sky130_fd_sc_hd__and2_4
XFILLER_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21424_ _15398_/Y _21285_/B VGND VGND VPWR VPWR _21424_/X sky130_fd_sc_hd__and2_4
XFILLER_136_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24212_ _23828_/CLK _16419_/X HRESETn VGND VGND VPWR VPWR _24212_/Q sky130_fd_sc_hd__dfrtp_4
X_25192_ _23085_/CLK _25192_/D HRESETn VGND VGND VPWR VPWR _25192_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25092__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24143_ _24113_/CLK _16591_/X HRESETn VGND VGND VPWR VPWR _24143_/Q sky130_fd_sc_hd__dfrtp_4
X_21355_ _17636_/X _21347_/X _21355_/C VGND VGND VPWR VPWR _21355_/X sky130_fd_sc_hd__or3_4
XFILLER_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20306_ _18614_/A _18614_/B VGND VGND VPWR VPWR _20306_/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25021__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24074_ _24079_/CLK _24074_/D HRESETn VGND VGND VPWR VPWR _16824_/A sky130_fd_sc_hd__dfrtp_4
X_21286_ _16551_/Y _21425_/B VGND VGND VPWR VPWR _21286_/X sky130_fd_sc_hd__and2_4
XFILLER_116_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23025_ _24189_/Q _23025_/B VGND VGND VPWR VPWR _23025_/Y sky130_fd_sc_hd__nor2_4
X_20237_ _23693_/Q _20251_/B _20236_/X VGND VGND VPWR VPWR _20237_/X sky130_fd_sc_hd__a21o_4
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15618__A3 _15505_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20168_ _20249_/A _20168_/B VGND VGND VPWR VPWR _20173_/A sky130_fd_sc_hd__and2_4
XFILLER_49_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11636__A _15801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19214__B1 _19170_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12990_ _12992_/A _12984_/B _12989_/Y VGND VGND VPWR VPWR _25012_/D sky130_fd_sc_hd__and3_4
X_20099_ _22106_/B _20098_/X _19597_/A _20098_/X VGND VGND VPWR VPWR _20099_/X sky130_fd_sc_hd__a2bb2o_4
X_24976_ _24980_/CLK _13389_/X HRESETn VGND VGND VPWR VPWR _24976_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11941_ _11940_/Y VGND VGND VPWR VPWR _11941_/X sky130_fd_sc_hd__buf_2
XFILLER_40_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23927_ _23469_/CLK _17940_/X HRESETn VGND VGND VPWR VPWR _23927_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16579__A1 _15799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14660_ _14657_/X _14659_/Y _15288_/A _14657_/X VGND VGND VPWR VPWR _24724_/D sky130_fd_sc_hd__a2bb2o_4
X_11872_ _25167_/Q _11871_/X _11869_/Y VGND VGND VPWR VPWR _11872_/X sky130_fd_sc_hd__o21a_4
X_23858_ _23767_/CLK _18296_/X HRESETn VGND VGND VPWR VPWR _23858_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_72_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13611_ _13611_/A VGND VGND VPWR VPWR _13611_/X sky130_fd_sc_hd__buf_2
X_22809_ _16492_/Y _20807_/X VGND VGND VPWR VPWR _22809_/X sky130_fd_sc_hd__and2_4
X_14591_ _14581_/A VGND VGND VPWR VPWR _18920_/A sky130_fd_sc_hd__buf_2
XFILLER_111_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23789_ _23789_/CLK _20692_/X HRESETn VGND VGND VPWR VPWR _23789_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22883__B _20807_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16330_ _24244_/Q VGND VGND VPWR VPWR _16330_/Y sky130_fd_sc_hd__inv_2
X_13542_ _23756_/Q _23755_/Q _23757_/Q _13541_/X VGND VGND VPWR VPWR _13543_/B sky130_fd_sc_hd__or4_4
XFILLER_38_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23956__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23060__A _20738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16261_ HWDATA[19] VGND VGND VPWR VPWR _16261_/X sky130_fd_sc_hd__buf_2
XFILLER_125_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13473_ _13473_/A VGND VGND VPWR VPWR _21257_/A sky130_fd_sc_hd__inv_2
X_18000_ _11630_/A VGND VGND VPWR VPWR _18000_/X sky130_fd_sc_hd__buf_2
X_15212_ _15108_/C _15216_/A VGND VGND VPWR VPWR _15213_/C sky130_fd_sc_hd__nand2_4
XFILLER_12_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12424_ _12424_/A _12424_/B VGND VGND VPWR VPWR _12424_/X sky130_fd_sc_hd__or2_4
XFILLER_12_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25109__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16192_ _16190_/Y _16191_/X _16100_/X _16191_/X VGND VGND VPWR VPWR _24300_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20835__B1 _20833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15143_ _15123_/A _15117_/C _14898_/Y VGND VGND VPWR VPWR _15143_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17993__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12355_ _22564_/A _12353_/Y _12403_/B _24472_/Q VGND VGND VPWR VPWR _12365_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12286_ _12267_/B VGND VGND VPWR VPWR _12287_/B sky130_fd_sc_hd__inv_2
X_15074_ _15067_/B _15071_/B VGND VGND VPWR VPWR _15075_/C sky130_fd_sc_hd__nand2_4
X_19951_ _19950_/Y _19948_/X _19421_/X _19948_/X VGND VGND VPWR VPWR _23149_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22588__B1 _22322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22404__A _22263_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14025_ _14618_/A _14037_/B VGND VGND VPWR VPWR _14025_/Y sky130_fd_sc_hd__nor2_4
X_18902_ _18897_/Y _18900_/X _18901_/X _18900_/X VGND VGND VPWR VPWR _18902_/X sky130_fd_sc_hd__a2bb2o_4
X_19882_ _19882_/A VGND VGND VPWR VPWR _22075_/B sky130_fd_sc_hd__inv_2
XANTENNA__16402__A _16426_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16267__B1 _16266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22123__B _21979_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18833_ _18832_/Y VGND VGND VPWR VPWR _18833_/X sky130_fd_sc_hd__buf_2
XFILLER_67_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24744__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18764_ _18763_/X VGND VGND VPWR VPWR _18764_/X sky130_fd_sc_hd__buf_2
X_15976_ _15975_/Y _15973_/X _15788_/X _15973_/X VGND VGND VPWR VPWR _24370_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20859__A _18263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17715_ _17889_/A _17715_/B _17715_/C VGND VGND VPWR VPWR _17724_/B sky130_fd_sc_hd__and3_4
X_14927_ _14925_/A _24257_/Q _15110_/B _14926_/Y VGND VGND VPWR VPWR _14927_/X sky130_fd_sc_hd__o22a_4
X_18695_ _18694_/Y _18692_/X _17202_/X _18692_/X VGND VGND VPWR VPWR _18695_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21563__B2 _21562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17646_ _17646_/A VGND VGND VPWR VPWR _21153_/A sky130_fd_sc_hd__buf_2
XFILLER_1_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14858_ _14880_/A _14859_/A _15022_/A _24145_/Q VGND VGND VPWR VPWR _14858_/X sky130_fd_sc_hd__a2bb2o_4
X_13809_ _13808_/X VGND VGND VPWR VPWR _13811_/C sky130_fd_sc_hd__inv_2
XANTENNA__13480__B _13480_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17577_ _17510_/B _17492_/X VGND VGND VPWR VPWR _17577_/X sky130_fd_sc_hd__or2_4
XFILLER_50_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14789_ _24710_/Q _14777_/Y _15059_/A _24097_/Q VGND VGND VPWR VPWR _14789_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20682__A1_N _20556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19316_ _23378_/Q VGND VGND VPWR VPWR _19316_/Y sky130_fd_sc_hd__inv_2
X_16528_ _16527_/Y _16523_/X _16100_/X _16523_/X VGND VGND VPWR VPWR _16528_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23697__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19247_ _21631_/B _19244_/X _11848_/X _19244_/X VGND VGND VPWR VPWR _19247_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16459_ _24196_/Q VGND VGND VPWR VPWR _16459_/Y sky130_fd_sc_hd__inv_2
X_19178_ _19177_/Y _19175_/X _19109_/X _19175_/X VGND VGND VPWR VPWR _23427_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22815__A1 _22195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22815__B2 _22198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11567__B1 _11566_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18129_ _23801_/Q _18112_/A _20886_/A _18125_/X VGND VGND VPWR VPWR _18129_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_8_104_0_HCLK clkbuf_7_52_0_HCLK/X VGND VGND VPWR VPWR _24412_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_117_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21140_ _21144_/A _21140_/B _21139_/X VGND VGND VPWR VPWR _21140_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_167_0_HCLK clkbuf_7_83_0_HCLK/X VGND VGND VPWR VPWR _25052_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_132_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21071_ _21066_/X _21070_/X _20782_/X VGND VGND VPWR VPWR _21071_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22001__A2_N _22259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12840__A _12951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16258__B1 _15855_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20022_ _23122_/Q VGND VGND VPWR VPWR _21605_/B sky130_fd_sc_hd__inv_2
XANTENNA__24485__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14808__B2 _24128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24830_ _24953_/CLK _24830_/D HRESETn VGND VGND VPWR VPWR _24830_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21872__B _15639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16273__A3 _15499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24414__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24761_ _24968_/CLK _14408_/X HRESETn VGND VGND VPWR VPWR _13438_/A sky130_fd_sc_hd__dfrtp_4
X_21973_ _24473_/Q _21543_/A VGND VGND VPWR VPWR _21973_/X sky130_fd_sc_hd__or2_4
XFILLER_132_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0_0_HCLK_A clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22751__B1 _20780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23712_ _23716_/CLK _23712_/D HRESETn VGND VGND VPWR VPWR _20499_/A sky130_fd_sc_hd__dfrtp_4
X_20924_ _21553_/A _20923_/X _20740_/A _13618_/A VGND VGND VPWR VPWR _20925_/A sky130_fd_sc_hd__o22a_4
XFILLER_15_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24692_ _24712_/CLK _24692_/D HRESETn VGND VGND VPWR VPWR _24692_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _21293_/B VGND VGND VPWR VPWR _22153_/B sky130_fd_sc_hd__buf_2
XFILLER_54_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23643_ _23641_/CLK scl_i_S4 HRESETn VGND VGND VPWR VPWR _23643_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22503__B1 _22351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16982__A _24046_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20786_ _20786_/A VGND VGND VPWR VPWR _20787_/B sky130_fd_sc_hd__buf_2
XPHY_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23574_ _23531_/CLK _23574_/D VGND VGND VPWR VPWR _17671_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22525_ _22129_/X _22524_/X _21994_/X _24411_/Q _21995_/X VGND VGND VPWR VPWR _22525_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12010__A1_N _12054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25202__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22456_ _22438_/X _22456_/B _22456_/C _22455_/Y VGND VGND VPWR VPWR _22456_/X sky130_fd_sc_hd__or4_4
XFILLER_108_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_63_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_63_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21407_ _21272_/X _21324_/X _21366_/X _21406_/X VGND VGND VPWR VPWR HRDATA[2] sky130_fd_sc_hd__or4_4
X_22387_ _22299_/A _22386_/X VGND VGND VPWR VPWR _22387_/X sky130_fd_sc_hd__and2_4
XFILLER_68_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25175_ _23100_/CLK _25175_/D HRESETn VGND VGND VPWR VPWR _19714_/A sky130_fd_sc_hd__dfrtp_4
X_12140_ _12133_/X _12140_/B _12137_/X _12139_/X VGND VGND VPWR VPWR _12140_/X sky130_fd_sc_hd__or4_4
XFILLER_68_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21338_ _21334_/X _21337_/X _17639_/X VGND VGND VPWR VPWR _21338_/X sky130_fd_sc_hd__o21a_4
X_24126_ _24101_/CLK _16618_/X HRESETn VGND VGND VPWR VPWR _24126_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12071_ _12071_/A VGND VGND VPWR VPWR _12178_/C sky130_fd_sc_hd__inv_2
X_21269_ _21269_/A _21710_/B VGND VGND VPWR VPWR _21269_/X sky130_fd_sc_hd__or2_4
XANTENNA__19435__B1 _19366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24057_ _24612_/CLK _24057_/D HRESETn VGND VGND VPWR VPWR _17021_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16249__B1 _24281_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23008_ _24498_/Q _23008_/B VGND VGND VPWR VPWR _23008_/X sky130_fd_sc_hd__or2_4
XANTENNA__17997__B1 _17205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15830_ _15830_/A VGND VGND VPWR VPWR _15830_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24155__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23055__A _23042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15761_ HWDATA[24] VGND VGND VPWR VPWR _15761_/X sky130_fd_sc_hd__buf_2
X_12973_ _21840_/A _12973_/B VGND VGND VPWR VPWR _12974_/B sky130_fd_sc_hd__or2_4
X_24959_ _24957_/CLK _24959_/D HRESETn VGND VGND VPWR VPWR _11653_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21545__A1 _11623_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17500_ _17581_/A _17494_/Y _17497_/X _17499_/X VGND VGND VPWR VPWR _17500_/X sky130_fd_sc_hd__or4_4
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21545__B2 _21544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14712_ _14874_/A VGND VGND VPWR VPWR _14712_/X sky130_fd_sc_hd__buf_2
XANTENNA__17053__A _17053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11924_ _11919_/A VGND VGND VPWR VPWR _11924_/X sky130_fd_sc_hd__buf_2
X_18480_ _18463_/A _18470_/B _18480_/C VGND VGND VPWR VPWR _18480_/X sky130_fd_sc_hd__and3_4
X_15692_ _15692_/A VGND VGND VPWR VPWR _16581_/A sky130_fd_sc_hd__buf_2
XFILLER_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17431_ _17411_/B _17431_/B _17428_/C VGND VGND VPWR VPWR _23983_/D sky130_fd_sc_hd__and3_4
X_14643_ _14643_/A VGND VGND VPWR VPWR _23685_/D sky130_fd_sc_hd__buf_2
XFILLER_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11855_ _11855_/A VGND VGND VPWR VPWR _19617_/A sky130_fd_sc_hd__buf_2
XFILLER_96_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17362_ _17362_/A _17362_/B _17361_/Y VGND VGND VPWR VPWR _17362_/X sky130_fd_sc_hd__and3_4
XFILLER_18_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14574_ _14565_/X VGND VGND VPWR VPWR _14574_/Y sky130_fd_sc_hd__inv_2
X_11786_ _11785_/X VGND VGND VPWR VPWR _11786_/Y sky130_fd_sc_hd__inv_2
X_19101_ _19114_/A VGND VGND VPWR VPWR _19101_/X sky130_fd_sc_hd__buf_2
XANTENNA__23790__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16313_ _16313_/A VGND VGND VPWR VPWR _16339_/A sky130_fd_sc_hd__buf_2
X_13525_ _13525_/A VGND VGND VPWR VPWR _13525_/Y sky130_fd_sc_hd__inv_2
X_17293_ _25218_/Q _17340_/A _11623_/Y _23982_/Q VGND VGND VPWR VPWR _17293_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16724__B2 _22376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19032_ _18068_/X VGND VGND VPWR VPWR _19799_/A sky130_fd_sc_hd__buf_2
X_16244_ _14920_/Y _16242_/X _16243_/X _16242_/X VGND VGND VPWR VPWR _16244_/X sky130_fd_sc_hd__a2bb2o_4
X_13456_ _13456_/A _14369_/B VGND VGND VPWR VPWR _13474_/B sky130_fd_sc_hd__and2_4
XANTENNA__11549__B1 _11548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12407_ _12406_/Y _12407_/B VGND VGND VPWR VPWR _12408_/D sky130_fd_sc_hd__or2_4
X_16175_ _16174_/Y _16170_/X _15777_/X _16170_/X VGND VGND VPWR VPWR _16175_/X sky130_fd_sc_hd__a2bb2o_4
X_13387_ _24853_/Q _13386_/X VGND VGND VPWR VPWR _13388_/B sky130_fd_sc_hd__or2_4
XANTENNA__24996__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20861__B _20861_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15126_ _15144_/A VGND VGND VPWR VPWR _15126_/X sky130_fd_sc_hd__buf_2
X_12338_ _25089_/Q VGND VGND VPWR VPWR _12412_/C sky130_fd_sc_hd__inv_2
XFILLER_86_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24925__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22134__A _25077_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15057_ _14982_/A VGND VGND VPWR VPWR _15057_/X sky130_fd_sc_hd__buf_2
X_19934_ _23155_/Q VGND VGND VPWR VPWR _21659_/B sky130_fd_sc_hd__inv_2
XANTENNA__19426__B1 _19424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12269_ _12103_/Y _12281_/B VGND VGND VPWR VPWR _12282_/B sky130_fd_sc_hd__or2_4
XFILLER_130_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14008_ _13925_/C _13950_/A VGND VGND VPWR VPWR _14008_/Y sky130_fd_sc_hd__nand2_4
XANTENNA_clkbuf_5_17_0_HCLK_A clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21973__A _24473_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19865_ _22071_/B _19864_/X _19815_/X _19864_/X VGND VGND VPWR VPWR _23182_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17988__B1 _15507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22981__B1 _17021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18816_ _13156_/B VGND VGND VPWR VPWR _18816_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19796_ _21235_/B _19793_/X _19462_/X _19793_/X VGND VGND VPWR VPWR _23208_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16660__B1 _15507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19729__B2 _19727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15959_ _22521_/A VGND VGND VPWR VPWR _15959_/Y sky130_fd_sc_hd__inv_2
X_18747_ _23579_/Q VGND VGND VPWR VPWR _18747_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22733__B1 _20782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13491__A _20883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18678_ HWDATA[3] VGND VGND VPWR VPWR _18678_/X sky130_fd_sc_hd__buf_2
XANTENNA__23878__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16412__B1 _15479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17629_ _23939_/Q _17629_/B VGND VGND VPWR VPWR _17630_/B sky130_fd_sc_hd__and2_4
XFILLER_91_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20640_ _23746_/Q _20635_/X _20644_/B VGND VGND VPWR VPWR _20640_/Y sky130_fd_sc_hd__a21oi_4
X_20571_ _23731_/Q _13529_/X _20570_/Y VGND VGND VPWR VPWR _20571_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16715__B2 _17615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22310_ _14047_/A _22307_/X _22308_/X _22310_/D VGND VGND VPWR VPWR _22310_/X sky130_fd_sc_hd__or4_4
X_23290_ _23112_/CLK _23290_/D VGND VGND VPWR VPWR _23290_/Q sky130_fd_sc_hd__dfxtp_4
X_22241_ _20909_/X _22239_/X _22240_/X _25200_/Q _21402_/X VGND VGND VPWR VPWR _22241_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21472__B1 _17639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22172_ _12328_/A _21565_/A VGND VGND VPWR VPWR _22172_/X sky130_fd_sc_hd__and2_4
XFILLER_118_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24666__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21123_ _21122_/X VGND VGND VPWR VPWR _21123_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22016__A2 _22014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16042__A _16042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22979__A _22979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21054_ _22249_/A VGND VGND VPWR VPWR _21710_/B sky130_fd_sc_hd__buf_2
XANTENNA__11712__B1 _11711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20005_ _13262_/B VGND VGND VPWR VPWR _20005_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_HCLK clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16651__B1 _15497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17994__A3 _17993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24813_ _24884_/CLK _24813_/D HRESETn VGND VGND VPWR VPWR _14234_/A sky130_fd_sc_hd__dfstp_4
XFILLER_132_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22724__B1 _14781_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24744_ _25052_/CLK _14537_/Y HRESETn VGND VGND VPWR VPWR _14528_/A sky130_fd_sc_hd__dfrtp_4
X_21956_ _14524_/B _21956_/B VGND VGND VPWR VPWR _21956_/X sky130_fd_sc_hd__or2_4
XANTENNA__16403__B1 _16243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _20833_/X _20906_/X VGND VGND VPWR VPWR _20907_/Y sky130_fd_sc_hd__nor2_4
XPHY_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24675_ _24676_/CLK _24675_/D HRESETn VGND VGND VPWR VPWR _24675_/Q sky130_fd_sc_hd__dfrtp_4
X_21887_ _21887_/A VGND VGND VPWR VPWR _21887_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _25190_/Q VGND VGND VPWR VPWR _11640_/Y sky130_fd_sc_hd__inv_2
XPHY_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23626_ _23624_/CLK _20708_/X HRESETn VGND VGND VPWR VPWR _20709_/A sky130_fd_sc_hd__dfstp_4
X_20838_ _15578_/B VGND VGND VPWR VPWR _20838_/X sky130_fd_sc_hd__buf_2
XPHY_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18156__B1 _16050_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22219__A _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11571_ _11568_/Y _11569_/X _11570_/X _11569_/X VGND VGND VPWR VPWR _25208_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16706__A1 _24367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23557_ _23133_/CLK _23557_/D VGND VGND VPWR VPWR _13061_/B sky130_fd_sc_hd__dfxtp_4
X_20769_ _20757_/X _20765_/X _22884_/B _20768_/X VGND VGND VPWR VPWR _20769_/X sky130_fd_sc_hd__a211o_4
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16706__B2 _17595_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13310_ _13102_/X _13308_/X _13310_/C VGND VGND VPWR VPWR _13310_/X sky130_fd_sc_hd__and3_4
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22508_ _24206_/Q _22574_/B _23023_/A VGND VGND VPWR VPWR _22508_/X sky130_fd_sc_hd__o21a_4
X_14290_ _24790_/Q VGND VGND VPWR VPWR _14290_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23488_ _23489_/CLK _23488_/D VGND VGND VPWR VPWR _19005_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__12464__B _12495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13241_ _13136_/A _13241_/B VGND VGND VPWR VPWR _13243_/B sky130_fd_sc_hd__or2_4
X_22439_ _16351_/Y _22439_/B VGND VGND VPWR VPWR _22439_/X sky130_fd_sc_hd__or2_4
XFILLER_13_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13172_ _13207_/A _13172_/B _13172_/C VGND VGND VPWR VPWR _13173_/C sky130_fd_sc_hd__or3_4
X_25158_ _25159_/CLK _11934_/X HRESETn VGND VGND VPWR VPWR _11933_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12594__A1_N _25054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12123_ _25119_/Q _12121_/Y _12180_/A _24550_/Q VGND VGND VPWR VPWR _12123_/X sky130_fd_sc_hd__a2bb2o_4
X_24109_ _24112_/CLK _16648_/X HRESETn VGND VGND VPWR VPWR _22502_/A sky130_fd_sc_hd__dfrtp_4
X_17980_ _17979_/X VGND VGND VPWR VPWR _17999_/A sky130_fd_sc_hd__inv_2
XANTENNA__24336__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_150_0_HCLK clkbuf_7_75_0_HCLK/X VGND VGND VPWR VPWR _25012_/CLK sky130_fd_sc_hd__clkbuf_1
X_25089_ _24488_/CLK _12476_/X HRESETn VGND VGND VPWR VPWR _25089_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20018__B2 _20015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12054_ _12054_/A _18111_/B VGND VGND VPWR VPWR _12054_/X sky130_fd_sc_hd__and2_4
X_16931_ _16834_/D _16927_/X VGND VGND VPWR VPWR _16931_/Y sky130_fd_sc_hd__nand2_4
XFILLER_77_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21793__A _21793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15791__A _15767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16862_ _16822_/A _16876_/A VGND VGND VPWR VPWR _16874_/B sky130_fd_sc_hd__or2_4
X_19650_ _21935_/B _19647_/X _19600_/X _19647_/X VGND VGND VPWR VPWR _19650_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22401__B _22265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15813_ _16222_/C _15729_/A _15810_/X _15812_/Y VGND VGND VPWR VPWR _15813_/X sky130_fd_sc_hd__a211o_4
X_18601_ _16320_/A _18438_/A _24242_/Q _18488_/A VGND VGND VPWR VPWR _18601_/X sky130_fd_sc_hd__a2bb2o_4
X_19581_ _19575_/Y VGND VGND VPWR VPWR _19581_/X sky130_fd_sc_hd__buf_2
X_16793_ _15849_/Y _16821_/A _15849_/Y _16821_/A VGND VGND VPWR VPWR _16793_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18532_ _18532_/A _18536_/A _18535_/A _18535_/B VGND VGND VPWR VPWR _18532_/X sky130_fd_sc_hd__or4_4
X_15744_ _16305_/A _15578_/X VGND VGND VPWR VPWR _15744_/X sky130_fd_sc_hd__or2_4
X_12956_ _12955_/X VGND VGND VPWR VPWR _12957_/B sky130_fd_sc_hd__inv_2
XFILLER_20_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23971__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11907_ _11905_/A _11884_/X _11906_/Y VGND VGND VPWR VPWR _20691_/A sky130_fd_sc_hd__o21a_4
X_18463_ _18463_/A _18461_/X _18462_/X VGND VGND VPWR VPWR _23840_/D sky130_fd_sc_hd__and3_4
XANTENNA__25195__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15675_ _15658_/X _15672_/X _15600_/X _24490_/Q _15661_/X VGND VGND VPWR VPWR _15675_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_2_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12887_ _12860_/Y _12894_/A _12963_/A _12886_/X VGND VGND VPWR VPWR _12890_/B sky130_fd_sc_hd__or4_4
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23900__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17414_ _17262_/Y _17423_/B VGND VGND VPWR VPWR _17421_/B sky130_fd_sc_hd__or2_4
XFILLER_60_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14626_ _14626_/A _14626_/B _24723_/Q VGND VGND VPWR VPWR _14627_/B sky130_fd_sc_hd__or3_4
XANTENNA__25124__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11838_ _19603_/A VGND VGND VPWR VPWR _11838_/Y sky130_fd_sc_hd__inv_2
X_18394_ _16418_/Y _23835_/Q _16448_/A _18425_/A VGND VGND VPWR VPWR _18394_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17345_ _17622_/B VGND VGND VPWR VPWR _17345_/X sky130_fd_sc_hd__buf_2
X_14557_ _17717_/A VGND VGND VPWR VPWR _17877_/A sky130_fd_sc_hd__buf_2
X_11769_ _11769_/A VGND VGND VPWR VPWR _17448_/A sky130_fd_sc_hd__inv_2
XANTENNA__19895__B1 _19828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16127__A _16127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13508_ _20468_/A _20469_/B _13508_/C _13508_/D VGND VGND VPWR VPWR _13509_/C sky130_fd_sc_hd__or4_4
X_17276_ _11583_/Y _17311_/A _11583_/Y _17311_/A VGND VGND VPWR VPWR _17277_/D sky130_fd_sc_hd__a2bb2o_4
X_14488_ _14487_/X VGND VGND VPWR VPWR _14488_/X sky130_fd_sc_hd__buf_2
X_19015_ _23485_/Q VGND VGND VPWR VPWR _21946_/B sky130_fd_sc_hd__inv_2
X_16227_ _14435_/B _16225_/Y _16003_/Y _16225_/Y VGND VGND VPWR VPWR _16227_/X sky130_fd_sc_hd__a2bb2o_4
X_13439_ _24933_/Q _13438_/A _13437_/Y _13438_/Y VGND VGND VPWR VPWR _13440_/D sky130_fd_sc_hd__o22a_4
XFILLER_31_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16158_ _16165_/A VGND VGND VPWR VPWR _16158_/X sky130_fd_sc_hd__buf_2
X_15109_ _24660_/Q VGND VGND VPWR VPWR _15109_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16089_ _24338_/Q VGND VGND VPWR VPWR _16089_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16476__A3 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24077__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19917_ _19917_/A VGND VGND VPWR VPWR _19917_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24006__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22954__B1 _20782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19848_ _21774_/B _19842_/X _19821_/X _19847_/X VGND VGND VPWR VPWR _23188_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16633__B1 HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19779_ _14493_/A _19779_/B _14548_/X _14549_/X VGND VGND VPWR VPWR _19780_/A sky130_fd_sc_hd__or4_4
X_21810_ _20967_/A _21808_/X _21810_/C VGND VGND VPWR VPWR _21810_/X sky130_fd_sc_hd__and3_4
X_22790_ _20819_/X _22788_/Y _22536_/X _22789_/X VGND VGND VPWR VPWR _22791_/A sky130_fd_sc_hd__o22a_4
XANTENNA__22965__C _22951_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21741_ _11938_/A _21300_/B _24777_/Q _23616_/Q _21088_/X VGND VGND VPWR VPWR _21741_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_25_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15739__A2 _15617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23641__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24460_ _24478_/CLK _24460_/D HRESETn VGND VGND VPWR VPWR _24460_/Q sky130_fd_sc_hd__dfrtp_4
X_21672_ _14471_/A _21672_/B _21671_/X VGND VGND VPWR VPWR _21672_/X sky130_fd_sc_hd__or3_4
Xclkbuf_4_13_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18354__A1_N _24211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23411_ _23411_/CLK _23411_/D VGND VGND VPWR VPWR _23411_/Q sky130_fd_sc_hd__dfxtp_4
X_20623_ _23742_/Q _20618_/X _20653_/A VGND VGND VPWR VPWR _20623_/Y sky130_fd_sc_hd__a21boi_4
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24391_ _24405_/CLK _15924_/X HRESETn VGND VGND VPWR VPWR _23002_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_20_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20554_ _20554_/A _20554_/B VGND VGND VPWR VPWR _20555_/A sky130_fd_sc_hd__or2_4
XFILLER_138_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23342_ _24748_/CLK _19419_/X VGND VGND VPWR VPWR _13032_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16694__A2_N _16692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20782__A _20782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24847__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15372__B1 _11590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20485_ _13509_/X VGND VGND VPWR VPWR _20517_/A sky130_fd_sc_hd__buf_2
X_23273_ _23249_/CLK _23273_/D VGND VGND VPWR VPWR _23273_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24026__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25012_ _25012_/CLK _25012_/D HRESETn VGND VGND VPWR VPWR _22133_/A sky130_fd_sc_hd__dfrtp_4
X_22224_ _22547_/A VGND VGND VPWR VPWR _22225_/A sky130_fd_sc_hd__buf_2
XANTENNA__21996__A1 _15322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22155_ _22155_/A _22155_/B _22155_/C VGND VGND VPWR VPWR _22155_/X sky130_fd_sc_hd__and3_4
XFILLER_105_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21106_ _20844_/B VGND VGND VPWR VPWR _21106_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_223_0_HCLK clkbuf_8_223_0_HCLK/A VGND VGND VPWR VPWR _24654_/CLK sky130_fd_sc_hd__clkbuf_1
X_22086_ _21626_/A _22084_/X _22085_/X VGND VGND VPWR VPWR _22086_/X sky130_fd_sc_hd__and3_4
XFILLER_120_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22502__A _22502_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17018__D _17017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22945__B1 _14740_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21037_ _21030_/X _21032_/X _21036_/X _24546_/Q _11530_/X VGND VGND VPWR VPWR _21038_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20420__B2 _20419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23729__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12810_ _22633_/A VGND VGND VPWR VPWR _12810_/Y sky130_fd_sc_hd__inv_2
X_13790_ _13779_/X _13789_/Y VGND VGND VPWR VPWR _13790_/X sky130_fd_sc_hd__or2_4
X_22988_ _16048_/A _22311_/A _22864_/X VGND VGND VPWR VPWR _22988_/X sky130_fd_sc_hd__o21a_4
XFILLER_28_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12741_ _12647_/B _12741_/B VGND VGND VPWR VPWR _12742_/B sky130_fd_sc_hd__or2_4
Xclkbuf_1_0_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_0_1_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_24727_ _23661_/CLK _14649_/X HRESETn VGND VGND VPWR VPWR _24727_/Q sky130_fd_sc_hd__dfrtp_4
X_21939_ _21227_/A _21939_/B VGND VGND VPWR VPWR _21939_/X sky130_fd_sc_hd__or2_4
X_15460_ _15689_/A VGND VGND VPWR VPWR _15460_/X sky130_fd_sc_hd__buf_2
X_12672_ _12578_/Y _12672_/B VGND VGND VPWR VPWR _12673_/C sky130_fd_sc_hd__or2_4
XFILLER_70_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24658_ _24662_/CLK _24658_/D HRESETn VGND VGND VPWR VPWR _24658_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _13413_/Y _14380_/B VGND VGND VPWR VPWR _14411_/Y sky130_fd_sc_hd__nand2_4
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _25194_/Q VGND VGND VPWR VPWR _11623_/Y sky130_fd_sc_hd__inv_2
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609_ _25050_/CLK _23609_/D VGND VGND VPWR VPWR _23609_/Q sky130_fd_sc_hd__dfxtp_4
X_15391_ _21888_/A _15387_/X _15390_/X _15387_/X VGND VGND VPWR VPWR _15391_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_54_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19877__B1 _19832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24589_ _23702_/CLK _24589_/D HRESETn VGND VGND VPWR VPWR _24589_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17130_ _17043_/B _17124_/X _17083_/X _17127_/B VGND VGND VPWR VPWR _17131_/A sky130_fd_sc_hd__a211o_4
XANTENNA__20487__A1 _13509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ _24774_/Q _14325_/A _24773_/Q _14319_/X VGND VGND VPWR VPWR _14342_/X sky130_fd_sc_hd__o22a_4
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11554_ _25213_/Q VGND VGND VPWR VPWR _11554_/Y sky130_fd_sc_hd__inv_2
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24588__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17061_ _17063_/B VGND VGND VPWR VPWR _17062_/B sky130_fd_sc_hd__inv_2
X_14273_ _14273_/A VGND VGND VPWR VPWR _14273_/X sky130_fd_sc_hd__buf_2
XANTENNA__24517__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16012_ _15438_/A _16006_/X _16008_/X _16224_/D VGND VGND VPWR VPWR _16012_/X sky130_fd_sc_hd__a211o_4
XFILLER_100_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13224_ _11710_/X _13208_/X _13223_/X _25000_/Q _13114_/X VGND VGND VPWR VPWR _13224_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__21436__B1 _13613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21300__B _21300_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_33_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_67_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_3_3_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13155_ _23893_/Q VGND VGND VPWR VPWR _13155_/X sky130_fd_sc_hd__buf_2
XANTENNA__17655__A2 _16222_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24170__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12106_ _12096_/X _12099_/X _12106_/C _12106_/D VGND VGND VPWR VPWR _12106_/X sky130_fd_sc_hd__or4_4
XFILLER_111_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13086_ _13171_/A _13083_/X _13085_/X VGND VGND VPWR VPWR _13087_/C sky130_fd_sc_hd__and3_4
X_17963_ _17899_/A _18895_/A VGND VGND VPWR VPWR _17963_/X sky130_fd_sc_hd__or2_4
XANTENNA__22936__B1 _22407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19702_ _19700_/Y _19701_/X _19614_/X _19701_/X VGND VGND VPWR VPWR _23241_/D sky130_fd_sc_hd__a2bb2o_4
X_12037_ _23798_/Q _12016_/X _12036_/Y VGND VGND VPWR VPWR _20698_/A sky130_fd_sc_hd__o21a_4
X_16914_ _16916_/B VGND VGND VPWR VPWR _16915_/B sky130_fd_sc_hd__inv_2
X_17894_ _17894_/A _17894_/B _17894_/C VGND VGND VPWR VPWR _17898_/B sky130_fd_sc_hd__and3_4
XANTENNA__16615__B1 _16291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19633_ _19633_/A VGND VGND VPWR VPWR _21469_/B sky130_fd_sc_hd__inv_2
XFILLER_38_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16845_ _16846_/A _16844_/Y VGND VGND VPWR VPWR _16845_/X sky130_fd_sc_hd__or2_4
XANTENNA__17225__B _11728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16091__B2 _16090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16776_ _16776_/A VGND VGND VPWR VPWR _16927_/A sky130_fd_sc_hd__inv_2
X_19564_ _23290_/Q VGND VGND VPWR VPWR _21477_/B sky130_fd_sc_hd__inv_2
XFILLER_59_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13988_ _13973_/X _13987_/Y _14234_/A _13938_/X VGND VGND VPWR VPWR _24885_/D sky130_fd_sc_hd__a2bb2o_4
X_15727_ _15712_/A _15720_/A VGND VGND VPWR VPWR _15728_/A sky130_fd_sc_hd__or2_4
X_18515_ _18515_/A _18515_/B VGND VGND VPWR VPWR _18518_/B sky130_fd_sc_hd__or2_4
X_12939_ _12880_/C _12937_/A VGND VGND VPWR VPWR _12939_/X sky130_fd_sc_hd__or2_4
X_19495_ _19493_/Y _19489_/X _19448_/X _19494_/X VGND VGND VPWR VPWR _19495_/X sky130_fd_sc_hd__a2bb2o_4
X_15658_ _15657_/X VGND VGND VPWR VPWR _15658_/X sky130_fd_sc_hd__buf_2
X_18446_ _18446_/A _18445_/X VGND VGND VPWR VPWR _18446_/X sky130_fd_sc_hd__or2_4
XFILLER_21_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14609_ _14609_/A _14683_/A _14681_/A _24718_/Q VGND VGND VPWR VPWR _14610_/B sky130_fd_sc_hd__or4_4
X_18377_ _18369_/X _18371_/X _18374_/X _18376_/X VGND VGND VPWR VPWR _18377_/X sky130_fd_sc_hd__or4_4
X_15589_ _15588_/Y VGND VGND VPWR VPWR _15593_/A sky130_fd_sc_hd__buf_2
X_17328_ _17353_/A _17305_/Y _17327_/X VGND VGND VPWR VPWR _17328_/X sky130_fd_sc_hd__or3_4
Xclkbuf_7_115_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_231_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24940__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17259_ _17252_/X _17259_/B _17259_/C _17258_/X VGND VGND VPWR VPWR _17259_/X sky130_fd_sc_hd__or4_4
XANTENNA__15354__B1 _11563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24258__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20270_ _24018_/Q _23657_/Q VGND VGND VPWR VPWR _23653_/D sky130_fd_sc_hd__and2_4
XANTENNA__11915__B1 _11913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11729__A _11728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22322__A _22322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23960_ _23949_/CLK _23960_/D HRESETn VGND VGND VPWR VPWR _23960_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23893__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12340__B1 _12412_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_53_0_HCLK clkbuf_8_53_0_HCLK/A VGND VGND VPWR VPWR _24944_/CLK sky130_fd_sc_hd__clkbuf_1
X_22911_ _21490_/X _22910_/X _22835_/X _25218_/Q _22840_/X VGND VGND VPWR VPWR _22911_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23891_ _24005_/CLK _18087_/X HRESETn VGND VGND VPWR VPWR _11732_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23822__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25046__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22842_ _22971_/A _22841_/X VGND VGND VPWR VPWR _22842_/X sky130_fd_sc_hd__and2_4
XFILLER_84_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20777__A _20749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22773_ _22769_/X _22773_/B _22773_/C _22772_/X VGND VGND VPWR VPWR _22773_/X sky130_fd_sc_hd__or4_4
XANTENNA__21902__B2 _20802_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17151__A _17129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24512_ _25005_/CLK _24512_/D HRESETn VGND VGND VPWR VPWR _24512_/Q sky130_fd_sc_hd__dfrtp_4
X_21724_ _13370_/Y _21707_/B _16462_/A _16041_/X VGND VGND VPWR VPWR _21724_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24443_ _24445_/CLK _24443_/D HRESETn VGND VGND VPWR VPWR _22420_/A sky130_fd_sc_hd__dfrtp_4
X_21655_ _21205_/A _21655_/B VGND VGND VPWR VPWR _21655_/X sky130_fd_sc_hd__or2_4
XFILLER_138_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20606_ _23738_/Q _20599_/A VGND VGND VPWR VPWR _20606_/X sky130_fd_sc_hd__or2_4
X_24374_ _24385_/CLK _15967_/X HRESETn VGND VGND VPWR VPWR _22436_/A sky130_fd_sc_hd__dfrtp_4
X_21586_ _11499_/A _21586_/B VGND VGND VPWR VPWR _21587_/C sky130_fd_sc_hd__or2_4
XANTENNA__24681__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23325_ _24748_/CLK _23325_/D VGND VGND VPWR VPWR _19470_/A sky130_fd_sc_hd__dfxtp_4
X_20537_ _20537_/A VGND VGND VPWR VPWR _23722_/D sky130_fd_sc_hd__inv_2
XFILLER_123_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24610__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20468_ _20468_/A VGND VGND VPWR VPWR _20468_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21120__B _13324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23256_ _23471_/CLK _23256_/D VGND VGND VPWR VPWR _19661_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_118_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22207_ _16041_/X VGND VGND VPWR VPWR _22931_/A sky130_fd_sc_hd__buf_2
XFILLER_134_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20399_ _20398_/X VGND VGND VPWR VPWR _20399_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14015__A _14015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23187_ _23493_/CLK _23187_/D VGND VGND VPWR VPWR _23187_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_134_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22138_ _22023_/X _22051_/X _22138_/C _22138_/D VGND VGND VPWR VPWR HRDATA[7] sky130_fd_sc_hd__or4_4
XANTENNA__13659__B1 _13658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14960_ _14960_/A VGND VGND VPWR VPWR _14960_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22069_ _21786_/A _19778_/Y VGND VGND VPWR VPWR _22070_/C sky130_fd_sc_hd__or2_4
XFILLER_121_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13911_ _13886_/A VGND VGND VPWR VPWR _13911_/X sky130_fd_sc_hd__buf_2
X_14891_ _14890_/Y VGND VGND VPWR VPWR _15138_/A sky130_fd_sc_hd__buf_2
XFILLER_134_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16630_ _14740_/Y _16629_/X HWDATA[29] _16629_/X VGND VGND VPWR VPWR _16630_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20848__A2_N _13614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13842_ _13811_/X _13822_/X _13833_/X _13841_/X VGND VGND VPWR VPWR _13842_/X sky130_fd_sc_hd__a211o_4
XFILLER_74_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16561_ _13614_/A VGND VGND VPWR VPWR _21590_/B sky130_fd_sc_hd__buf_2
XFILLER_16_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23063__A _20741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13773_ _13730_/X _24637_/Q _13773_/C _13773_/D VGND VGND VPWR VPWR _13774_/B sky130_fd_sc_hd__or4_4
X_15512_ _12111_/Y _15509_/X _15511_/X _15509_/X VGND VGND VPWR VPWR _24554_/D sky130_fd_sc_hd__a2bb2o_4
X_18300_ _18300_/A _18327_/A _18167_/Y _18299_/X VGND VGND VPWR VPWR _18301_/B sky130_fd_sc_hd__or4_4
X_12724_ _12644_/D _12700_/B _12674_/X _12722_/B VGND VGND VPWR VPWR _12725_/A sky130_fd_sc_hd__a211o_4
X_19280_ _19279_/Y _19274_/X _19232_/X _19260_/X VGND VGND VPWR VPWR _19280_/X sky130_fd_sc_hd__a2bb2o_4
X_16492_ _16492_/A VGND VGND VPWR VPWR _16492_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24769__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18231_ _18258_/A _18222_/D VGND VGND VPWR VPWR _18231_/X sky130_fd_sc_hd__or2_4
X_15443_ _14436_/B _15443_/B VGND VGND VPWR VPWR _15443_/X sky130_fd_sc_hd__or2_4
X_12655_ _12550_/X _12571_/Y _12642_/X _12654_/X VGND VGND VPWR VPWR _12655_/X sky130_fd_sc_hd__or4_4
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11606_ _25198_/Q VGND VGND VPWR VPWR _11606_/Y sky130_fd_sc_hd__inv_2
X_18162_ _16078_/A _23863_/Q _16078_/Y _18279_/A VGND VGND VPWR VPWR _18163_/D sky130_fd_sc_hd__o22a_4
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15374_ _15358_/X VGND VGND VPWR VPWR _15374_/X sky130_fd_sc_hd__buf_2
XFILLER_30_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12586_ _12584_/A _12585_/A _12584_/Y _12585_/Y VGND VGND VPWR VPWR _12586_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16128__A2 _16135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21121__A2 _11952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17113_ _17101_/A _17108_/X _17112_/X VGND VGND VPWR VPWR _17113_/X sky130_fd_sc_hd__and3_4
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14325_ _14325_/A VGND VGND VPWR VPWR _14325_/X sky130_fd_sc_hd__buf_2
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11537_ _11537_/A VGND VGND VPWR VPWR _11537_/X sky130_fd_sc_hd__buf_2
X_18093_ _18093_/A _18092_/X VGND VGND VPWR VPWR _18093_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15336__B1 _11540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24351__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17044_ _17124_/B _17044_/B VGND VGND VPWR VPWR _17044_/X sky130_fd_sc_hd__or2_4
XFILLER_7_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21409__B1 _24548_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14256_ _14255_/Y _14253_/X _14209_/X _14253_/X VGND VGND VPWR VPWR _14256_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13207_ _13207_/A _13207_/B _13207_/C VGND VGND VPWR VPWR _13208_/C sky130_fd_sc_hd__or3_4
X_14187_ _14174_/Y _14186_/X _11975_/A _14180_/X VGND VGND VPWR VPWR _24827_/D sky130_fd_sc_hd__o22a_4
XFILLER_124_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13138_ _13090_/X _13138_/B _13138_/C VGND VGND VPWR VPWR _13138_/X sky130_fd_sc_hd__and3_4
X_18995_ _23492_/Q VGND VGND VPWR VPWR _21763_/B sky130_fd_sc_hd__inv_2
XFILLER_39_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13069_ _13078_/A VGND VGND VPWR VPWR _13169_/A sky130_fd_sc_hd__buf_2
X_17946_ _17914_/A _17944_/X _17946_/C VGND VGND VPWR VPWR _17947_/C sky130_fd_sc_hd__and3_4
XFILLER_65_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16081__A1_N _16080_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21981__A _22629_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17877_ _17877_/A _23449_/Q VGND VGND VPWR VPWR _17877_/X sky130_fd_sc_hd__or2_4
XFILLER_93_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17261__B1 _11524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19616_ _19616_/A VGND VGND VPWR VPWR _21146_/B sky130_fd_sc_hd__inv_2
XFILLER_26_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16828_ _16760_/Y _16800_/Y _16885_/A VGND VGND VPWR VPWR _16840_/A sky130_fd_sc_hd__or3_4
XFILLER_38_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19547_ _21328_/B _19546_/X _11857_/X _19546_/X VGND VGND VPWR VPWR _19547_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16759_ _24405_/Q _16834_/D _15841_/Y _24085_/Q VGND VGND VPWR VPWR _16759_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19478_ _19477_/Y _19473_/X _19360_/X _19473_/X VGND VGND VPWR VPWR _23322_/D sky130_fd_sc_hd__a2bb2o_4
X_18429_ _23825_/Q VGND VGND VPWR VPWR _18515_/A sky130_fd_sc_hd__inv_2
XANTENNA__24439__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13004__A _12925_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21440_ _12004_/Y _13357_/X _18122_/Y _21083_/X VGND VGND VPWR VPWR _21440_/X sky130_fd_sc_hd__o22a_4
XFILLER_124_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22317__A _22263_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21371_ _21371_/A _19938_/Y VGND VGND VPWR VPWR _21372_/C sky130_fd_sc_hd__or2_4
XANTENNA__24092__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22860__A2 _22859_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20322_ _24805_/Q _18624_/A VGND VGND VPWR VPWR _20322_/X sky130_fd_sc_hd__or2_4
X_23110_ _23293_/CLK _20053_/X VGND VGND VPWR VPWR _23110_/Q sky130_fd_sc_hd__dfxtp_4
X_24090_ _24088_/CLK _24090_/D HRESETn VGND VGND VPWR VPWR _16846_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_31_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20253_ _23659_/Q _23770_/Q _23772_/Q _23771_/Q VGND VGND VPWR VPWR _20254_/D sky130_fd_sc_hd__or4_4
XFILLER_116_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23041_ _23041_/A _20881_/A VGND VGND VPWR VPWR _23041_/X sky130_fd_sc_hd__and2_4
XANTENNA__21875__B _20885_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20623__A1 _23742_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20184_ _14206_/A _20182_/X _20178_/A _20183_/X VGND VGND VPWR VPWR _20184_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_130_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24992_ _24841_/CLK _24992_/D HRESETn VGND VGND VPWR VPWR _24992_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21891__A _24822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23943_ _23972_/CLK _17621_/X HRESETn VGND VGND VPWR VPWR _16720_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12864__B2 _24432_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23874_ _24641_/CLK _18236_/X HRESETn VGND VGND VPWR VPWR _18234_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20139__B1 _19421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22825_ _22637_/X _22822_/Y _22601_/X _22824_/X VGND VGND VPWR VPWR _22825_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21115__B _21867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22756_ _22348_/X _22749_/X _22751_/X _22585_/X _22755_/Y VGND VGND VPWR VPWR _22756_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24862__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14942__A2_N _24269_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21707_ _21707_/A _21707_/B VGND VGND VPWR VPWR _21707_/X sky130_fd_sc_hd__or2_4
XFILLER_90_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22687_ _22665_/Y _22687_/B _22687_/C _22686_/X VGND VGND VPWR VPWR HRDATA[20] sky130_fd_sc_hd__or4_4
X_12440_ _12417_/A _12438_/A VGND VGND VPWR VPWR _12440_/X sky130_fd_sc_hd__or2_4
XFILLER_100_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24426_ _24425_/CLK _15829_/X HRESETn VGND VGND VPWR VPWR _24426_/Q sky130_fd_sc_hd__dfrtp_4
X_21638_ _21638_/A VGND VGND VPWR VPWR _21638_/X sky130_fd_sc_hd__buf_2
XANTENNA__24109__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21131__A _17629_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12371_ _22564_/A VGND VGND VPWR VPWR _12412_/B sky130_fd_sc_hd__inv_2
X_24357_ _25183_/CLK _24357_/D HRESETn VGND VGND VPWR VPWR _16014_/B sky130_fd_sc_hd__dfrtp_4
X_21569_ _21569_/A _21569_/B _21568_/X VGND VGND VPWR VPWR _21569_/X sky130_fd_sc_hd__and3_4
XANTENNA__12753__A _12749_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14957__A2_N _24259_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14110_ _13391_/B _11916_/X _13388_/B VGND VGND VPWR VPWR _14110_/X sky130_fd_sc_hd__or3_4
XANTENNA__20862__A1 _16294_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23308_ _23308_/CLK _19517_/X VGND VGND VPWR VPWR _23308_/Q sky130_fd_sc_hd__dfxtp_4
X_15090_ _15087_/A _15093_/B VGND VGND VPWR VPWR _15090_/Y sky130_fd_sc_hd__nand2_4
X_24288_ _23353_/CLK _24288_/D HRESETn VGND VGND VPWR VPWR _15435_/A sky130_fd_sc_hd__dfrtp_4
X_14041_ _14041_/A VGND VGND VPWR VPWR _20719_/A sky130_fd_sc_hd__inv_2
X_23239_ _23356_/CLK _23239_/D VGND VGND VPWR VPWR _23239_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13287__C _13287_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16879__B _17067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23058__A _20736_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23744__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17800_ _17903_/A _18949_/A VGND VGND VPWR VPWR _17800_/X sky130_fd_sc_hd__or2_4
XFILLER_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15992_ _13632_/A VGND VGND VPWR VPWR _15992_/X sky130_fd_sc_hd__buf_2
X_18780_ _17956_/B VGND VGND VPWR VPWR _18780_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12304__B1 _12508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14943_ _14935_/X _14943_/B _14943_/C _14943_/D VGND VGND VPWR VPWR _14943_/X sky130_fd_sc_hd__or4_4
X_17731_ _17780_/A _17731_/B _17731_/C VGND VGND VPWR VPWR _17738_/B sky130_fd_sc_hd__and3_4
XFILLER_48_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14874_ _14874_/A VGND VGND VPWR VPWR _14874_/Y sky130_fd_sc_hd__inv_2
X_17662_ _17662_/A _17662_/B _17655_/X VGND VGND VPWR VPWR _17663_/A sky130_fd_sc_hd__or3_4
XFILLER_75_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22119__A1 _22116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22119__B2 _22118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19401_ _13146_/B VGND VGND VPWR VPWR _19401_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13825_ _24906_/Q VGND VGND VPWR VPWR _13825_/X sky130_fd_sc_hd__buf_2
X_16613_ _14835_/Y _16610_/X _16546_/X _16610_/X VGND VGND VPWR VPWR _16613_/X sky130_fd_sc_hd__a2bb2o_4
X_17593_ _17603_/A _17591_/X _17593_/C VGND VGND VPWR VPWR _23953_/D sky130_fd_sc_hd__and3_4
X_16544_ _16544_/A VGND VGND VPWR VPWR _16544_/Y sky130_fd_sc_hd__inv_2
X_19332_ _19331_/Y _19328_/X _19308_/X _19328_/X VGND VGND VPWR VPWR _23373_/D sky130_fd_sc_hd__a2bb2o_4
X_13756_ _13769_/D VGND VGND VPWR VPWR _13782_/B sky130_fd_sc_hd__buf_2
XFILLER_95_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12707_ _12707_/A VGND VGND VPWR VPWR _12707_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17207__A2_N _17198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16475_ _16475_/A _16475_/B VGND VGND VPWR VPWR _16475_/X sky130_fd_sc_hd__or2_4
X_19263_ _19263_/A VGND VGND VPWR VPWR _19263_/Y sky130_fd_sc_hd__inv_2
X_13687_ _13686_/X VGND VGND VPWR VPWR _13687_/X sky130_fd_sc_hd__buf_2
XANTENNA__24532__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15426_ _20861_/B VGND VGND VPWR VPWR _15426_/X sky130_fd_sc_hd__buf_2
X_18214_ _23849_/Q VGND VGND VPWR VPWR _18214_/Y sky130_fd_sc_hd__inv_2
X_12638_ _24462_/Q VGND VGND VPWR VPWR _12638_/Y sky130_fd_sc_hd__inv_2
X_19194_ _19193_/Y _19191_/X _19149_/X _19191_/X VGND VGND VPWR VPWR _19194_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19299__B2 _19296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21041__A _20751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15357_ _15357_/A VGND VGND VPWR VPWR _22587_/A sky130_fd_sc_hd__inv_2
X_18145_ _18145_/A _18145_/B _18145_/C _18145_/D VGND VGND VPWR VPWR _18164_/B sky130_fd_sc_hd__or4_4
X_12569_ _24510_/Q VGND VGND VPWR VPWR _12569_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14780__B2 _14779_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16135__A _16134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14308_ _20164_/A VGND VGND VPWR VPWR _20185_/A sky130_fd_sc_hd__buf_2
X_18076_ _18075_/X VGND VGND VPWR VPWR _18690_/B sky130_fd_sc_hd__buf_2
XFILLER_116_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15288_ _15288_/A VGND VGND VPWR VPWR _15288_/Y sky130_fd_sc_hd__inv_2
X_17027_ _17027_/A VGND VGND VPWR VPWR _17133_/A sky130_fd_sc_hd__inv_2
X_14239_ _24812_/Q VGND VGND VPWR VPWR _14239_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23037__A2_N _21491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18978_ _18977_/Y _18975_/X _18953_/X _18975_/X VGND VGND VPWR VPWR _18978_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14296__B1 _14209_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17929_ _17929_/A _17929_/B _17929_/C VGND VGND VPWR VPWR _17929_/X sky130_fd_sc_hd__and3_4
XFILLER_117_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20908__A2 _22497_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20940_ _20902_/X VGND VGND VPWR VPWR _20940_/X sky130_fd_sc_hd__buf_2
XFILLER_94_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20871_ _20701_/A _21638_/A _20269_/B _21088_/A VGND VGND VPWR VPWR _20871_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_82_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15796__B1 _15393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_127_0_HCLK clkbuf_7_63_0_HCLK/X VGND VGND VPWR VPWR _23762_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__11742__A _11741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22610_ _22610_/A VGND VGND VPWR VPWR _22610_/X sky130_fd_sc_hd__buf_2
XPHY_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23590_ _23457_/CLK _23590_/D VGND VGND VPWR VPWR _17701_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_81_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_6_0_HCLK_A clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22541_ _21540_/X _22538_/X _20839_/X _22540_/X VGND VGND VPWR VPWR _22541_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24273__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22472_ _22306_/A _22462_/X _22465_/X _22471_/X VGND VGND VPWR VPWR _22472_/X sky130_fd_sc_hd__or4_4
XFILLER_37_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24202__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24211_ _24262_/CLK _24211_/D HRESETn VGND VGND VPWR VPWR _24211_/Q sky130_fd_sc_hd__dfrtp_4
X_21423_ _20566_/Y _22279_/A _20429_/Y _22610_/A VGND VGND VPWR VPWR _21423_/X sky130_fd_sc_hd__o22a_4
X_25191_ _24405_/CLK _11639_/X HRESETn VGND VGND VPWR VPWR _25191_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21886__A _20926_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24142_ _24145_/CLK _16592_/X HRESETn VGND VGND VPWR VPWR _24142_/Q sky130_fd_sc_hd__dfrtp_4
X_21354_ _21350_/X _21353_/X _21172_/X VGND VGND VPWR VPWR _21355_/C sky130_fd_sc_hd__o21a_4
X_20305_ _20305_/A VGND VGND VPWR VPWR _23635_/D sky130_fd_sc_hd__inv_2
XANTENNA__15884__A _24404_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24073_ _24079_/CLK _24073_/D HRESETn VGND VGND VPWR VPWR _16825_/A sky130_fd_sc_hd__dfrtp_4
X_21285_ _21285_/A _21285_/B VGND VGND VPWR VPWR _21285_/X sky130_fd_sc_hd__and2_4
XFILLER_11_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23024_ _23726_/Q _22285_/X _23758_/Q _22531_/X VGND VGND VPWR VPWR _23024_/Y sky130_fd_sc_hd__a22oi_4
X_20236_ _24822_/Q _14309_/X _20234_/X _20192_/X _20235_/X VGND VGND VPWR VPWR _20236_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_81_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20167_ _20167_/A VGND VGND VPWR VPWR _20168_/B sky130_fd_sc_hd__inv_2
XANTENNA__25061__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14826__A2 _24155_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18017__A2 _15657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20098_ _20110_/A VGND VGND VPWR VPWR _20098_/X sky130_fd_sc_hd__buf_2
X_24975_ _24980_/CLK _24975_/D HRESETn VGND VGND VPWR VPWR SCLK_S2 sky130_fd_sc_hd__dfstp_4
XANTENNA__12837__B2 _22385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11940_ _20847_/A VGND VGND VPWR VPWR _11940_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17604__A _17595_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23926_ _23442_/CLK _23926_/D HRESETn VGND VGND VPWR VPWR _23926_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_23_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18973__B1 _18880_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21126__A _13334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_86_0_HCLK clkbuf_7_87_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_86_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_11871_ _11871_/A _11871_/B _11871_/C _11871_/D VGND VGND VPWR VPWR _11871_/X sky130_fd_sc_hd__and4_4
X_23857_ _23767_/CLK _23857_/D HRESETn VGND VGND VPWR VPWR _18209_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_73_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13610_ _16301_/A _13609_/X VGND VGND VPWR VPWR _13611_/A sky130_fd_sc_hd__or2_4
X_22808_ _24247_/Q _21553_/X _20780_/X _22807_/X VGND VGND VPWR VPWR _22808_/X sky130_fd_sc_hd__a211o_4
X_14590_ _14589_/B VGND VGND VPWR VPWR _14592_/B sky130_fd_sc_hd__inv_2
XFILLER_38_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23788_ _24984_/CLK _23788_/D HRESETn VGND VGND VPWR VPWR _11905_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_41_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18725__B1 _18679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13541_ _13540_/X VGND VGND VPWR VPWR _13541_/X sky130_fd_sc_hd__buf_2
XFILLER_125_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22739_ _16501_/Y _21576_/X _15347_/Y _22452_/X VGND VGND VPWR VPWR _22739_/X sky130_fd_sc_hd__o22a_4
X_16260_ _14958_/Y _16257_/X _16259_/X _16257_/X VGND VGND VPWR VPWR _16260_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13472_ _13461_/X VGND VGND VPWR VPWR _19946_/B sky130_fd_sc_hd__buf_2
X_15211_ _15192_/A _15211_/B _15210_/Y VGND VGND VPWR VPWR _24658_/D sky130_fd_sc_hd__and3_4
XANTENNA__14896__A2_N _24271_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12423_ _12423_/A _12399_/A VGND VGND VPWR VPWR _12424_/B sky130_fd_sc_hd__and2_4
X_24409_ _24412_/CLK _24409_/D HRESETn VGND VGND VPWR VPWR _24409_/Q sky130_fd_sc_hd__dfrtp_4
X_16191_ _16196_/A VGND VGND VPWR VPWR _16191_/X sky130_fd_sc_hd__buf_2
XFILLER_138_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19150__B1 _19149_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23996__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15142_ _15154_/A _15140_/X _15141_/X VGND VGND VPWR VPWR _24677_/D sky130_fd_sc_hd__and3_4
XANTENNA__20835__A1 _16305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12354_ _25075_/Q VGND VGND VPWR VPWR _12403_/B sky130_fd_sc_hd__inv_2
XFILLER_127_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23925__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15073_ _14743_/X _15075_/B _15072_/Y VGND VGND VPWR VPWR _24691_/D sky130_fd_sc_hd__o21a_4
X_19950_ _23149_/Q VGND VGND VPWR VPWR _19950_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25149__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12285_ _12281_/B _12285_/B _12300_/C VGND VGND VPWR VPWR _12285_/X sky130_fd_sc_hd__and3_4
XANTENNA__15711__B1 _20808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22588__A1 _22011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14024_ _20396_/A VGND VGND VPWR VPWR _14618_/A sky130_fd_sc_hd__inv_2
X_18901_ _18763_/X VGND VGND VPWR VPWR _18901_/X sky130_fd_sc_hd__buf_2
XFILLER_106_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19881_ _21008_/B _19876_/X _19859_/X _19876_/A VGND VGND VPWR VPWR _19881_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18832_ _18832_/A VGND VGND VPWR VPWR _18832_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14278__B1 _14221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18763_ HWDATA[7] VGND VGND VPWR VPWR _18763_/X sky130_fd_sc_hd__buf_2
XFILLER_23_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15975_ _22239_/A VGND VGND VPWR VPWR _15975_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17216__B1 _16617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20859__B _20861_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17714_ _17853_/A _17714_/B VGND VGND VPWR VPWR _17715_/C sky130_fd_sc_hd__or2_4
X_14926_ _24257_/Q VGND VGND VPWR VPWR _14926_/Y sky130_fd_sc_hd__inv_2
X_18694_ _23597_/Q VGND VGND VPWR VPWR _18694_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24784__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21563__A2 _21561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17645_ _23938_/Q VGND VGND VPWR VPWR _17646_/A sky130_fd_sc_hd__inv_2
XANTENNA__15778__B1 _15777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14857_ _14697_/Y _24156_/Q _14697_/Y _24156_/Q VGND VGND VPWR VPWR _14857_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24713__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14849__A2_N _14836_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15034__A _15034_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13808_ _13808_/A VGND VGND VPWR VPWR _13808_/X sky130_fd_sc_hd__buf_2
X_14788_ _14977_/C _24123_/Q _14977_/C _24123_/Q VGND VGND VPWR VPWR _14788_/X sky130_fd_sc_hd__a2bb2o_4
X_17576_ _17575_/X VGND VGND VPWR VPWR _23956_/D sky130_fd_sc_hd__inv_2
XFILLER_63_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20118__A3 _13663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19315_ _19314_/Y _19312_/X _19221_/X _19312_/X VGND VGND VPWR VPWR _23379_/D sky130_fd_sc_hd__a2bb2o_4
X_13739_ _13745_/A _13725_/Y _13735_/X _13737_/Y _13738_/X VGND VGND VPWR VPWR _13739_/X
+ sky130_fd_sc_hd__a32o_4
X_16527_ _16527_/A VGND VGND VPWR VPWR _16527_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19246_ _19246_/A VGND VGND VPWR VPWR _21631_/B sky130_fd_sc_hd__inv_2
XFILLER_34_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16458_ _16457_/Y _16452_/X _16369_/X _16452_/X VGND VGND VPWR VPWR _16458_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15409_ _21113_/B VGND VGND VPWR VPWR _22024_/B sky130_fd_sc_hd__buf_2
X_16389_ _16389_/A VGND VGND VPWR VPWR _16389_/Y sky130_fd_sc_hd__inv_2
X_19177_ _19177_/A VGND VGND VPWR VPWR _19177_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14753__B2 _24098_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18128_ _18127_/Y _18125_/X _20886_/A _18125_/X VGND VGND VPWR VPWR _23879_/D sky130_fd_sc_hd__a2bb2o_4
X_18059_ _23903_/Q _17634_/A _19530_/A _17634_/Y VGND VGND VPWR VPWR _18059_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18080__A _18080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22314__B _22314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21070_ _21067_/Y _22322_/A _13526_/A _21069_/X VGND VGND VPWR VPWR _21070_/X sky130_fd_sc_hd__a2bb2o_4
X_20021_ _21809_/B _20015_/X _19717_/X _20020_/X VGND VGND VPWR VPWR _23123_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14269__B1 _14228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17207__B1 _17205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22200__B1 _22167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21533__A1_N _21400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24760_ _24968_/CLK _24760_/D HRESETn VGND VGND VPWR VPWR _13435_/A sky130_fd_sc_hd__dfrtp_4
X_21972_ _20783_/X VGND VGND VPWR VPWR _21972_/X sky130_fd_sc_hd__buf_2
XANTENNA__22687__D _22686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17271__A1_N _25207_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23711_ _24604_/CLK _23711_/D HRESETn VGND VGND VPWR VPWR _20499_/C sky130_fd_sc_hd__dfrtp_4
X_20923_ _21179_/A _20922_/X _13519_/A _12062_/X VGND VGND VPWR VPWR _20923_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15769__B1 _15350_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24691_ _24264_/CLK _24691_/D HRESETn VGND VGND VPWR VPWR _24691_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24454__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23642_ _23648_/CLK _20330_/Y HRESETn VGND VGND VPWR VPWR _23642_/Q sky130_fd_sc_hd__dfrtp_4
X_20854_ _21432_/A VGND VGND VPWR VPWR _22444_/B sky130_fd_sc_hd__buf_2
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20785__A _13614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22503__A1 _24271_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15784__A3 _16093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23573_ _23531_/CLK _18767_/X VGND VGND VPWR VPWR _17743_/B sky130_fd_sc_hd__dfxtp_4
X_20785_ _13614_/X VGND VGND VPWR VPWR _20786_/A sky130_fd_sc_hd__buf_2
XPHY_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22524_ _24305_/Q _22524_/B VGND VGND VPWR VPWR _22524_/X sky130_fd_sc_hd__or2_4
XFILLER_50_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16194__B1 _15788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19297__A2_N _19296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22455_ _22455_/A VGND VGND VPWR VPWR _22455_/Y sky130_fd_sc_hd__inv_2
X_21406_ _21397_/Y _21405_/Y _21793_/A VGND VGND VPWR VPWR _21406_/X sky130_fd_sc_hd__o21a_4
XFILLER_109_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25174_ _23388_/CLK _25174_/D HRESETn VGND VGND VPWR VPWR _11837_/A sky130_fd_sc_hd__dfrtp_4
X_22386_ _21248_/X _22385_/X _22240_/X _24515_/Q _20780_/A VGND VGND VPWR VPWR _22386_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22505__A _22505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22019__B1 _16608_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24125_ _24104_/CLK _16619_/X HRESETn VGND VGND VPWR VPWR _24125_/Q sky130_fd_sc_hd__dfrtp_4
X_21337_ _21147_/A _21337_/B _21337_/C VGND VGND VPWR VPWR _21337_/X sky130_fd_sc_hd__and3_4
XFILLER_135_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12070_ _20889_/A _12067_/Y _11643_/X _12067_/Y VGND VGND VPWR VPWR _25134_/D sky130_fd_sc_hd__a2bb2o_4
X_24056_ _24055_/CLK _17064_/X HRESETn VGND VGND VPWR VPWR _24056_/Q sky130_fd_sc_hd__dfrtp_4
X_21268_ _21268_/A VGND VGND VPWR VPWR _21268_/Y sky130_fd_sc_hd__inv_2
X_23007_ _23006_/X VGND VGND VPWR VPWR _23007_/Y sky130_fd_sc_hd__inv_2
X_20219_ _20254_/A _20241_/A VGND VGND VPWR VPWR _20232_/C sky130_fd_sc_hd__and2_4
XFILLER_133_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19814__A _19831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21199_ _21234_/A VGND VGND VPWR VPWR _21393_/A sky130_fd_sc_hd__buf_2
XFILLER_133_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19199__B1 _19109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15760_ _15748_/X _15740_/X _15596_/X _24454_/Q _15746_/X VGND VGND VPWR VPWR _15760_/X
+ sky130_fd_sc_hd__a32o_4
X_12972_ _12972_/A _12972_/B VGND VGND VPWR VPWR _12973_/B sky130_fd_sc_hd__or2_4
X_24958_ _24957_/CLK _24958_/D HRESETn VGND VGND VPWR VPWR _24958_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21545__A2 _11986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18946__B1 _18901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11923_ _11923_/A VGND VGND VPWR VPWR _21707_/A sky130_fd_sc_hd__inv_2
X_14711_ _24692_/Q _14709_/Y _14880_/A _22857_/A VGND VGND VPWR VPWR _14719_/B sky130_fd_sc_hd__a2bb2o_4
X_15691_ _15684_/X _15689_/X _15505_/X _22373_/A _15685_/X VGND VGND VPWR VPWR _24479_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_2_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23909_ _24944_/CLK _23909_/D HRESETn VGND VGND VPWR VPWR _18005_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24195__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24889_ _23774_/CLK _13976_/X HRESETn VGND VGND VPWR VPWR _13928_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14642_ _14636_/X _14641_/X _24729_/Q _14636_/X VGND VGND VPWR VPWR _14642_/X sky130_fd_sc_hd__a2bb2o_4
X_17430_ _17430_/A _17430_/B VGND VGND VPWR VPWR _17431_/B sky130_fd_sc_hd__or2_4
X_11854_ _11851_/Y _11852_/X _11853_/X _11852_/X VGND VGND VPWR VPWR _25171_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24124__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22768__A2_N _22765_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_110_0_HCLK clkbuf_7_55_0_HCLK/X VGND VGND VPWR VPWR _24161_/CLK sky130_fd_sc_hd__clkbuf_1
X_14573_ _14573_/A _14555_/X VGND VGND VPWR VPWR _14573_/X sky130_fd_sc_hd__and2_4
X_17361_ _17255_/Y _17358_/B VGND VGND VPWR VPWR _17361_/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11785_ _11769_/A _11773_/C _11802_/C _11803_/C VGND VGND VPWR VPWR _11785_/X sky130_fd_sc_hd__a211o_4
XANTENNA__20505__B1 _20446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14693__A pwm_S6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_173_0_HCLK clkbuf_7_86_0_HCLK/X VGND VGND VPWR VPWR _25106_/CLK sky130_fd_sc_hd__clkbuf_1
X_19100_ _19100_/A _19100_/B VGND VGND VPWR VPWR _19114_/A sky130_fd_sc_hd__nor2_4
X_13524_ _23748_/Q _13524_/B _23749_/Q _13524_/D VGND VGND VPWR VPWR _20653_/B sky130_fd_sc_hd__or4_4
X_16312_ _16312_/A VGND VGND VPWR VPWR _16312_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17292_ _11496_/Y _24008_/Q _11496_/Y _24008_/Q VGND VGND VPWR VPWR _17295_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16185__B1 _15369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16243_ HWDATA[29] VGND VGND VPWR VPWR _16243_/X sky130_fd_sc_hd__buf_2
X_19031_ _13022_/B VGND VGND VPWR VPWR _19031_/Y sky130_fd_sc_hd__inv_2
X_13455_ _13454_/X VGND VGND VPWR VPWR _14369_/B sky130_fd_sc_hd__inv_2
XFILLER_103_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15932__B1 _15837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12406_ _25080_/Q VGND VGND VPWR VPWR _12406_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13102__A _13299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16174_ _24306_/Q VGND VGND VPWR VPWR _16174_/Y sky130_fd_sc_hd__inv_2
X_13386_ _14107_/A _14108_/A _11917_/D _24852_/Q VGND VGND VPWR VPWR _13386_/X sky130_fd_sc_hd__and4_4
XFILLER_86_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15125_ _15125_/A _15125_/B VGND VGND VPWR VPWR _15125_/X sky130_fd_sc_hd__or2_4
X_12337_ _12327_/X _12337_/B _12337_/C _12336_/X VGND VGND VPWR VPWR _12337_/X sky130_fd_sc_hd__or4_4
XFILLER_138_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22134__B _20814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15056_ _15055_/X VGND VGND VPWR VPWR _15056_/Y sky130_fd_sc_hd__inv_2
X_19933_ _21766_/B _19927_/X _19448_/A _19932_/X VGND VGND VPWR VPWR _23156_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12268_ _12157_/Y _12283_/B VGND VGND VPWR VPWR _12281_/B sky130_fd_sc_hd__or2_4
X_14007_ _14007_/A VGND VGND VPWR VPWR _24881_/D sky130_fd_sc_hd__inv_2
XFILLER_96_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19864_ _19876_/A VGND VGND VPWR VPWR _19864_/X sky130_fd_sc_hd__buf_2
XANTENNA__21973__B _21543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12199_ _12198_/X VGND VGND VPWR VPWR _12200_/B sky130_fd_sc_hd__inv_2
XFILLER_110_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24965__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18815_ _18813_/Y _18809_/X _18744_/X _18814_/X VGND VGND VPWR VPWR _18815_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19795_ _19795_/A VGND VGND VPWR VPWR _21235_/B sky130_fd_sc_hd__inv_2
XFILLER_7_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18746_ _18742_/Y _18736_/X _18744_/X _18745_/X VGND VGND VPWR VPWR _23580_/D sky130_fd_sc_hd__a2bb2o_4
X_15958_ _15957_/Y _15953_/X _15777_/X _15953_/X VGND VGND VPWR VPWR _15958_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22733__A1 _24417_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14788__A2_N _24123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14909_ _24658_/Q VGND VGND VPWR VPWR _15108_/B sky130_fd_sc_hd__inv_2
XFILLER_23_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18677_ _23602_/Q VGND VGND VPWR VPWR _18677_/Y sky130_fd_sc_hd__inv_2
X_15889_ _15889_/A VGND VGND VPWR VPWR _15889_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17628_ _23938_/Q VGND VGND VPWR VPWR _17629_/B sky130_fd_sc_hd__buf_2
XFILLER_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14711__A2_N _14709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17559_ _16708_/Y _17564_/B _16748_/X VGND VGND VPWR VPWR _17559_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__12985__B1 _12896_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20570_ _13531_/B VGND VGND VPWR VPWR _20570_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23847__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19229_ _23408_/Q VGND VGND VPWR VPWR _21252_/A sky130_fd_sc_hd__inv_2
XFILLER_108_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22240_ _22646_/A VGND VGND VPWR VPWR _22240_/X sky130_fd_sc_hd__buf_2
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22171_ _13506_/D _22170_/X VGND VGND VPWR VPWR _22175_/B sky130_fd_sc_hd__and2_4
XFILLER_69_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21122_ _20885_/X _21117_/X _21119_/X _21120_/X _21121_/X VGND VGND VPWR VPWR _21122_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_28_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21053_ _21590_/B VGND VGND VPWR VPWR _22249_/A sky130_fd_sc_hd__buf_2
XANTENNA__22421__B1 _20801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20004_ _20002_/Y _20003_/X _19808_/X _20003_/X VGND VGND VPWR VPWR _20004_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24635__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24812_ _24884_/CLK _14240_/X HRESETn VGND VGND VPWR VPWR _24812_/Q sky130_fd_sc_hd__dfstp_4
X_24743_ _25052_/CLK _24743_/D HRESETn VGND VGND VPWR VPWR _14441_/A sky130_fd_sc_hd__dfrtp_4
X_21955_ _21376_/A _21955_/B _21955_/C VGND VGND VPWR VPWR _21955_/X sky130_fd_sc_hd__and3_4
XFILLER_76_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20906_ _20823_/X _20905_/X _23910_/Q _12063_/X VGND VGND VPWR VPWR _20906_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17600__B1 _16748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24674_ _24674_/CLK _24674_/D HRESETn VGND VGND VPWR VPWR _24674_/Q sky130_fd_sc_hd__dfrtp_4
X_21886_ _20926_/X VGND VGND VPWR VPWR _21886_/X sky130_fd_sc_hd__buf_2
XFILLER_42_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15105__C _14950_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23625_ _23624_/CLK _20706_/X HRESETn VGND VGND VPWR VPWR _20710_/B sky130_fd_sc_hd__dfstp_4
X_20837_ _20800_/X VGND VGND VPWR VPWR _20837_/X sky130_fd_sc_hd__buf_2
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14965__B2 _14936_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19353__B1 _19308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ HWDATA[18] VGND VGND VPWR VPWR _11570_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_246_0_HCLK clkbuf_8_247_0_HCLK/A VGND VGND VPWR VPWR _24712_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23556_ _23133_/CLK _18815_/X VGND VGND VPWR VPWR _23556_/Q sky130_fd_sc_hd__dfxtp_4
X_20768_ _16218_/Y _22445_/B VGND VGND VPWR VPWR _20768_/X sky130_fd_sc_hd__and2_4
XANTENNA__14851__A1_N _24706_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22507_ _16345_/A _22505_/X _20821_/X _22506_/X VGND VGND VPWR VPWR _22507_/X sky130_fd_sc_hd__a211o_4
XFILLER_35_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23487_ _23489_/CLK _19008_/X VGND VGND VPWR VPWR _23487_/Q sky130_fd_sc_hd__dfxtp_4
X_20699_ _12043_/X _20697_/B VGND VGND VPWR VPWR _23799_/D sky130_fd_sc_hd__and2_4
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13240_ _13155_/X _13232_/X _13240_/C VGND VGND VPWR VPWR _13240_/X sky130_fd_sc_hd__and3_4
X_22438_ _22438_/A _22434_/X _22437_/X VGND VGND VPWR VPWR _22438_/X sky130_fd_sc_hd__and3_4
XFILLER_87_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13171_ _13171_/A _13168_/X _13171_/C VGND VGND VPWR VPWR _13172_/C sky130_fd_sc_hd__and3_4
X_25157_ _25159_/CLK _11935_/X HRESETn VGND VGND VPWR VPWR _20880_/A sky130_fd_sc_hd__dfrtp_4
X_22369_ _21432_/A VGND VGND VPWR VPWR _22369_/X sky130_fd_sc_hd__buf_2
XFILLER_2_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12122_ _12122_/A VGND VGND VPWR VPWR _12180_/A sky130_fd_sc_hd__inv_2
X_24108_ _24113_/CLK _16651_/X HRESETn VGND VGND VPWR VPWR _16649_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_2_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25088_ _25091_/CLK _25088_/D HRESETn VGND VGND VPWR VPWR _25088_/Q sky130_fd_sc_hd__dfrtp_4
X_12053_ _12053_/A VGND VGND VPWR VPWR _12053_/Y sky130_fd_sc_hd__inv_2
X_16930_ _16834_/C _16932_/B _16929_/Y VGND VGND VPWR VPWR _24070_/D sky130_fd_sc_hd__o21a_4
X_24039_ _24612_/CLK _17131_/Y HRESETn VGND VGND VPWR VPWR _24039_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_5_9_0_HCLK_A clkbuf_4_4_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16861_ _16920_/A _16840_/B _16802_/Y _16840_/A VGND VGND VPWR VPWR _16876_/A sky130_fd_sc_hd__or4_4
XFILLER_81_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24376__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18600_ _16320_/Y _23839_/Q _16336_/Y _23833_/Q VGND VGND VPWR VPWR _18602_/C sky130_fd_sc_hd__a2bb2o_4
X_15812_ _15811_/X VGND VGND VPWR VPWR _15812_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17064__A _17052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19580_ _23284_/Q VGND VGND VPWR VPWR _21786_/B sky130_fd_sc_hd__inv_2
X_16792_ _15875_/Y _16829_/A _15875_/Y _16829_/A VGND VGND VPWR VPWR _16792_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24305__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22715__B2 _22657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18531_ _18543_/A _18543_/B VGND VGND VPWR VPWR _18535_/B sky130_fd_sc_hd__or2_4
XFILLER_93_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12955_ _12833_/X _12955_/B VGND VGND VPWR VPWR _12955_/X sky130_fd_sc_hd__or2_4
X_15743_ HWDATA[31] VGND VGND VPWR VPWR _15743_/X sky130_fd_sc_hd__buf_2
XFILLER_92_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11906_ _11905_/X VGND VGND VPWR VPWR _11906_/Y sky130_fd_sc_hd__inv_2
X_18462_ _18462_/A _18460_/A VGND VGND VPWR VPWR _18462_/X sky130_fd_sc_hd__or2_4
X_12886_ _12779_/Y _12885_/X VGND VGND VPWR VPWR _12886_/X sky130_fd_sc_hd__or2_4
X_15674_ _12332_/Y _15669_/X _11552_/X _15669_/X VGND VGND VPWR VPWR _15674_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_56_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_56_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17413_ _17413_/A _17413_/B VGND VGND VPWR VPWR _17423_/B sky130_fd_sc_hd__or2_4
X_11837_ _11837_/A VGND VGND VPWR VPWR _19603_/A sky130_fd_sc_hd__buf_2
X_14625_ _14625_/A _14625_/B _24721_/Q VGND VGND VPWR VPWR _14626_/B sky130_fd_sc_hd__or3_4
X_18393_ _18387_/X _18389_/X _18390_/X _18392_/X VGND VGND VPWR VPWR _18407_/B sky130_fd_sc_hd__or4_4
XANTENNA__12936__A _12854_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18147__A1 _16075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19344__B1 _19207_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11840__A _11830_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14556_ _14555_/X VGND VGND VPWR VPWR _14561_/A sky130_fd_sc_hd__inv_2
X_17344_ _17362_/A _17344_/B _17343_/X VGND VGND VPWR VPWR _17344_/X sky130_fd_sc_hd__and3_4
X_11768_ _21188_/A _11763_/X _11767_/X VGND VGND VPWR VPWR _11768_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_105_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23940__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ _23705_/Q _13506_/X VGND VGND VPWR VPWR _20469_/B sky130_fd_sc_hd__or2_4
XANTENNA__13445__A1_N _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14487_ _14486_/X VGND VGND VPWR VPWR _14487_/X sky130_fd_sc_hd__buf_2
X_17275_ _11592_/Y _23990_/Q _11592_/Y _23990_/Q VGND VGND VPWR VPWR _17277_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15905__B1 _15801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14708__B2 _22502_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25164__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11699_ _11706_/A _11696_/X _11701_/C _11698_/X VGND VGND VPWR VPWR _25189_/D sky130_fd_sc_hd__o22a_4
X_19014_ _19009_/Y _19013_/X _15541_/X _19013_/X VGND VGND VPWR VPWR _23486_/D sky130_fd_sc_hd__a2bb2o_4
X_13438_ _13438_/A VGND VGND VPWR VPWR _13438_/Y sky130_fd_sc_hd__inv_2
X_16226_ _16003_/Y _16225_/Y _14431_/A _16225_/Y VGND VGND VPWR VPWR _24288_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22145__A _21570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14870__B _15087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16157_ _24313_/Q VGND VGND VPWR VPWR _16157_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21454__A1 _12389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13369_ _21884_/A _13366_/X _11616_/X _13366_/X VGND VGND VPWR VPWR _24983_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15108_ _15208_/A _15108_/B _15108_/C _14969_/Y VGND VGND VPWR VPWR _15108_/X sky130_fd_sc_hd__or4_4
X_16088_ _22479_/A _16084_/X _16087_/X _16084_/X VGND VGND VPWR VPWR _24339_/D sky130_fd_sc_hd__a2bb2o_4
X_15039_ _15018_/X _15034_/X _15039_/C VGND VGND VPWR VPWR _24699_/D sky130_fd_sc_hd__and3_4
X_19916_ _21518_/B _19911_/X _19828_/X _19911_/X VGND VGND VPWR VPWR _19916_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15982__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24625__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22954__A1 _24424_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19847_ _19841_/X VGND VGND VPWR VPWR _19847_/X sky130_fd_sc_hd__buf_2
XFILLER_25_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19778_ _23214_/Q VGND VGND VPWR VPWR _19778_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24046__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18729_ _18728_/Y _18724_/X _18685_/X _18724_/X VGND VGND VPWR VPWR _18729_/X sky130_fd_sc_hd__a2bb2o_4
X_21740_ _14234_/Y _20818_/A _24805_/Q _20866_/A VGND VGND VPWR VPWR _21740_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16397__B1 _15320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22965__D _22964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15739__A3 _15735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21224__A _21224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21671_ _21665_/X _21670_/X _14440_/X VGND VGND VPWR VPWR _21671_/X sky130_fd_sc_hd__o21a_4
XFILLER_12_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14947__B2 _24278_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19335__B1 _19311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16318__A _24249_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23410_ _23411_/CLK _23410_/D VGND VGND VPWR VPWR _19223_/A sky130_fd_sc_hd__dfxtp_4
X_20622_ _13537_/C VGND VGND VPWR VPWR _20653_/A sky130_fd_sc_hd__buf_2
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24390_ _24590_/CLK _15926_/X HRESETn VGND VGND VPWR VPWR _24390_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23681__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23341_ _24748_/CLK _19422_/X VGND VGND VPWR VPWR _23341_/Q sky130_fd_sc_hd__dfxtp_4
X_20553_ _20552_/X VGND VGND VPWR VPWR _20553_/X sky130_fd_sc_hd__buf_2
XANTENNA__21693__B2 _15430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19629__A _19636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_13_0_HCLK clkbuf_7_6_0_HCLK/X VGND VGND VPWR VPWR _23336_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22770__A1_N _12415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_76_0_HCLK clkbuf_8_77_0_HCLK/A VGND VGND VPWR VPWR _24984_/CLK sky130_fd_sc_hd__clkbuf_1
X_23272_ _23249_/CLK _23272_/D VGND VGND VPWR VPWR _19616_/A sky130_fd_sc_hd__dfxtp_4
X_20484_ _20511_/A VGND VGND VPWR VPWR _20484_/X sky130_fd_sc_hd__buf_2
XANTENNA__15911__A3 _15735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25011_ _24435_/CLK _12992_/X HRESETn VGND VGND VPWR VPWR _25011_/Q sky130_fd_sc_hd__dfrtp_4
X_22223_ _22223_/A VGND VGND VPWR VPWR _22730_/A sky130_fd_sc_hd__buf_2
XANTENNA__21445__B2 _15426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17149__A _17129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24887__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24913__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22154_ _16107_/Y _22154_/B VGND VGND VPWR VPWR _22155_/C sky130_fd_sc_hd__or2_4
XFILLER_121_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24816__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21105_ _17614_/A _11516_/B _25006_/Q _21050_/Y VGND VGND VPWR VPWR _21105_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15892__A _15892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22085_ _21617_/A _22085_/B VGND VGND VPWR VPWR _22085_/X sky130_fd_sc_hd__or2_4
XANTENNA__22945__A1 _16400_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21036_ _22646_/A VGND VGND VPWR VPWR _21036_/X sky130_fd_sc_hd__buf_2
XFILLER_87_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22987_ _16398_/A _23020_/B VGND VGND VPWR VPWR _22990_/B sky130_fd_sc_hd__or2_4
XFILLER_103_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12740_ _12647_/C _12739_/X VGND VGND VPWR VPWR _12741_/B sky130_fd_sc_hd__or2_4
X_21938_ _21339_/A _21930_/X _21937_/X VGND VGND VPWR VPWR _21938_/X sky130_fd_sc_hd__and3_4
XFILLER_27_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16388__B1 _16219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20184__A1 _14206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24726_ _23661_/CLK _14652_/X HRESETn VGND VGND VPWR VPWR _24726_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_128_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23769__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12671_ _25066_/Q _12671_/B VGND VGND VPWR VPWR _12673_/B sky130_fd_sc_hd__or2_4
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24657_ _24662_/CLK _24657_/D HRESETn VGND VGND VPWR VPWR _14915_/A sky130_fd_sc_hd__dfrtp_4
X_21869_ _21866_/Y _20819_/X _22584_/A _21868_/X VGND VGND VPWR VPWR _21870_/B sky130_fd_sc_hd__o22a_4
XANTENNA__14938__B2 _14937_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18129__A1 _23801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16228__A _16228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14382_/B _14399_/X _14409_/Y _14403_/X _13435_/A VGND VGND VPWR VPWR _24760_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _11618_/Y _11610_/X _11620_/X _11621_/X VGND VGND VPWR VPWR _11622_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23608_ _25050_/CLK _18660_/X VGND VGND VPWR VPWR _23608_/Q sky130_fd_sc_hd__dfxtp_4
X_15390_ _16373_/A VGND VGND VPWR VPWR _15390_/X sky130_fd_sc_hd__buf_2
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17337__C1 _17336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24588_ _24013_/CLK _15397_/X HRESETn VGND VGND VPWR VPWR _15395_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ _14335_/X _14340_/X _14297_/A _14331_/X VGND VGND VPWR VPWR _14341_/X sky130_fd_sc_hd__o22a_4
XFILLER_11_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ _11550_/Y _11551_/X _11552_/X _11551_/X VGND VGND VPWR VPWR _11553_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20487__A2 _20481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23539_ _23133_/CLK _18862_/X VGND VGND VPWR VPWR _13157_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17060_ _17067_/A _17046_/X _17022_/B _17070_/A VGND VGND VPWR VPWR _17063_/B sky130_fd_sc_hd__or4_4
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14272_ _14272_/A VGND VGND VPWR VPWR _14272_/Y sky130_fd_sc_hd__inv_2
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16011_ _16011_/A VGND VGND VPWR VPWR _16224_/D sky130_fd_sc_hd__inv_2
X_13223_ _13113_/A _13215_/X _13222_/X VGND VGND VPWR VPWR _13223_/X sky130_fd_sc_hd__and3_4
XANTENNA__21436__A1 _21300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25209_ _25214_/CLK _25209_/D HRESETn VGND VGND VPWR VPWR _11565_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_137_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13154_ _13057_/X _13153_/X _25001_/Q _13116_/X VGND VGND VPWR VPWR _25001_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24557__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12105_ _25109_/Q _24552_/Q _12103_/Y _12104_/Y VGND VGND VPWR VPWR _12106_/D sky130_fd_sc_hd__o22a_4
X_13085_ _13085_/A _13085_/B VGND VGND VPWR VPWR _13085_/X sky130_fd_sc_hd__or2_4
X_17962_ _17815_/A _17962_/B _17961_/X VGND VGND VPWR VPWR _17970_/B sky130_fd_sc_hd__or3_4
XANTENNA__22936__A1 _13337_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19701_ _19688_/Y VGND VGND VPWR VPWR _19701_/X sky130_fd_sc_hd__buf_2
X_12036_ _12035_/X VGND VGND VPWR VPWR _12036_/Y sky130_fd_sc_hd__inv_2
X_16913_ _16839_/B _16912_/X VGND VGND VPWR VPWR _16916_/B sky130_fd_sc_hd__or2_4
X_17893_ _17782_/A _23561_/Q VGND VGND VPWR VPWR _17894_/C sky130_fd_sc_hd__or2_4
X_19632_ _21615_/B _19629_/X _19607_/X _19629_/X VGND VGND VPWR VPWR _23267_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16844_ _16816_/Y _16843_/X VGND VGND VPWR VPWR _16844_/Y sky130_fd_sc_hd__nor2_4
XFILLER_120_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19563_ _21624_/B _19560_/X _11848_/X _19560_/X VGND VGND VPWR VPWR _23291_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16775_ _24424_/Q _16774_/A _15832_/Y _16774_/Y VGND VGND VPWR VPWR _16775_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13987_ _13986_/X VGND VGND VPWR VPWR _13987_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18514_ _18468_/C _18485_/D VGND VGND VPWR VPWR _18515_/B sky130_fd_sc_hd__or2_4
XFILLER_80_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15726_ _15726_/A VGND VGND VPWR VPWR _15726_/Y sky130_fd_sc_hd__inv_2
X_12938_ _22712_/A _12937_/Y VGND VGND VPWR VPWR _12938_/X sky130_fd_sc_hd__or2_4
X_19494_ _19488_/Y VGND VGND VPWR VPWR _19494_/X sky130_fd_sc_hd__buf_2
XFILLER_20_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18445_ _18468_/C _18448_/A VGND VGND VPWR VPWR _18445_/X sky130_fd_sc_hd__and2_4
X_15657_ _15692_/A VGND VGND VPWR VPWR _15657_/X sky130_fd_sc_hd__buf_2
X_12869_ _22921_/A VGND VGND VPWR VPWR _12899_/C sky130_fd_sc_hd__inv_2
XFILLER_61_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19317__B1 _19201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16139__A2_N _16138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11570__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14608_ _24729_/Q VGND VGND VPWR VPWR _14608_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21979__A _21848_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18376_ _24192_/Q _23815_/Q _16469_/Y _18552_/A VGND VGND VPWR VPWR _18376_/X sky130_fd_sc_hd__o22a_4
X_15588_ _15584_/A VGND VGND VPWR VPWR _15588_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20883__A _20883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17327_ _17306_/Y _17255_/Y _17308_/X _17327_/D VGND VGND VPWR VPWR _17327_/X sky130_fd_sc_hd__or4_4
X_14539_ _24742_/Q VGND VGND VPWR VPWR _14539_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22872__B1 _22407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17258_ _25197_/Q _17257_/A _11609_/Y _17317_/C VGND VGND VPWR VPWR _17258_/X sky130_fd_sc_hd__o22a_4
XFILLER_31_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21427__A1 _13335_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13365__B1 _11607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16209_ _16207_/Y _16203_/X _15992_/X _16208_/X VGND VGND VPWR VPWR _16209_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13399__A1_N SSn_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17189_ _17171_/X _17185_/X _24025_/Q _24026_/Q _17188_/X VGND VGND VPWR VPWR _17189_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24980__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16303__B1 _16219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24298__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24227__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18056__B1 _21363_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20938__B1 _22011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11662__A2_N _23917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22910_ _22910_/A _22834_/B VGND VGND VPWR VPWR _22910_/X sky130_fd_sc_hd__or2_4
X_23890_ _23990_/CLK _23890_/D HRESETn VGND VGND VPWR VPWR _23890_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22841_ _21490_/X _22838_/X _22839_/X _25216_/Q _22840_/X VGND VGND VPWR VPWR _22841_/X
+ sky130_fd_sc_hd__a32o_4
X_22772_ _20520_/Y _22610_/X _20656_/A _22657_/X VGND VGND VPWR VPWR _22772_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23862__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24511_ _25005_/CLK _24511_/D HRESETn VGND VGND VPWR VPWR _12582_/A sky130_fd_sc_hd__dfrtp_4
X_21723_ _21722_/X VGND VGND VPWR VPWR _21723_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25086__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22992__B _22992_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24442_ _24445_/CLK _24442_/D HRESETn VGND VGND VPWR VPWR _22385_/A sky130_fd_sc_hd__dfrtp_4
X_21654_ _21238_/A _21654_/B VGND VGND VPWR VPWR _21654_/X sky130_fd_sc_hd__or2_4
XANTENNA__25015__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20793__A _22953_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20605_ _23738_/Q VGND VGND VPWR VPWR _20605_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15887__A _24403_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24373_ _24385_/CLK _15969_/X HRESETn VGND VGND VPWR VPWR _24373_/Q sky130_fd_sc_hd__dfrtp_4
X_21585_ _11890_/Y _22840_/A _21581_/X _22006_/B VGND VGND VPWR VPWR _21585_/X sky130_fd_sc_hd__a211o_4
XANTENNA__18263__A _18263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23324_ _24748_/CLK _19474_/X VGND VGND VPWR VPWR _23324_/Q sky130_fd_sc_hd__dfxtp_4
X_20536_ _22884_/A _20416_/A _20511_/A _20535_/X VGND VGND VPWR VPWR _20537_/A sky130_fd_sc_hd__o22a_4
XANTENNA__12159__B2 _24548_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13356__B1 _13330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23255_ _23356_/CLK _23255_/D VGND VGND VPWR VPWR _19663_/A sky130_fd_sc_hd__dfxtp_4
X_20467_ _20461_/X _20463_/Y _24594_/Q _20466_/X VGND VGND VPWR VPWR _20467_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22206_ _11985_/Y _11954_/X _14744_/A _22879_/A VGND VGND VPWR VPWR _22206_/X sky130_fd_sc_hd__a2bb2o_4
X_23186_ _23179_/CLK _23186_/D VGND VGND VPWR VPWR _23186_/Q sky130_fd_sc_hd__dfxtp_4
X_20398_ _14639_/Y _20343_/Y _20357_/X _20397_/Y VGND VGND VPWR VPWR _20398_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24650__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22137_ _22306_/A _22120_/X _22125_/X _22132_/X _22136_/X VGND VGND VPWR VPWR _22138_/D
+ sky130_fd_sc_hd__o41a_4
XFILLER_121_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20641__A2 _20552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16511__A _16499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22232__B _22265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22068_ _22055_/X _19967_/Y VGND VGND VPWR VPWR _22068_/X sky130_fd_sc_hd__or2_4
XFILLER_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11655__A _21871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13910_ _13806_/X _13908_/X _13905_/X _13845_/A _13903_/X VGND VGND VPWR VPWR _24903_/D
+ sky130_fd_sc_hd__a32o_4
X_21019_ _21019_/A VGND VGND VPWR VPWR _21020_/B sky130_fd_sc_hd__inv_2
XANTENNA__19822__A _19831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14890_ _24675_/Q VGND VGND VPWR VPWR _14890_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13841_ _13837_/X _13840_/Y _13837_/X _13840_/Y VGND VGND VPWR VPWR _13841_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_121_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_243_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13772_ _24649_/Q _13732_/A _13728_/X VGND VGND VPWR VPWR _13773_/C sky130_fd_sc_hd__or3_4
X_16560_ _15430_/X _16276_/X _16558_/X _15099_/A _16559_/X VGND VGND VPWR VPWR _24157_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_43_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21354__B1 _21172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15511_ HWDATA[9] VGND VGND VPWR VPWR _15511_/X sky130_fd_sc_hd__buf_2
XFILLER_128_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12723_ _12716_/A _12710_/D _12722_/X VGND VGND VPWR VPWR _25052_/D sky130_fd_sc_hd__and3_4
X_24709_ _24676_/CLK _24709_/D HRESETn VGND VGND VPWR VPWR _14997_/A sky130_fd_sc_hd__dfrtp_4
X_16491_ _16490_/Y _16486_/X _16153_/X _16486_/X VGND VGND VPWR VPWR _16491_/X sky130_fd_sc_hd__a2bb2o_4
X_18230_ _18229_/X VGND VGND VPWR VPWR _18230_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12654_ _12646_/X _12653_/X VGND VGND VPWR VPWR _12654_/X sky130_fd_sc_hd__or2_4
X_15442_ RsRx_S0 _15440_/A _15452_/B VGND VGND VPWR VPWR _15443_/B sky130_fd_sc_hd__o21a_4
XFILLER_128_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ _11603_/Y _11599_/X _11604_/X _11599_/X VGND VGND VPWR VPWR _11605_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18161_ _23863_/Q VGND VGND VPWR VPWR _18279_/A sky130_fd_sc_hd__inv_2
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _12585_/A VGND VGND VPWR VPWR _12585_/Y sky130_fd_sc_hd__inv_2
X_15373_ _15373_/A VGND VGND VPWR VPWR _22344_/A sky130_fd_sc_hd__inv_2
XFILLER_128_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17112_ _16992_/A _17112_/B VGND VGND VPWR VPWR _17112_/X sky130_fd_sc_hd__or2_4
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11536_ HWDATA[28] VGND VGND VPWR VPWR _11536_/X sky130_fd_sc_hd__buf_2
X_14324_ _23650_/Q VGND VGND VPWR VPWR _14325_/A sky130_fd_sc_hd__buf_2
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18092_ _18091_/Y _11766_/Y _21644_/A _17226_/X VGND VGND VPWR VPWR _18092_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16533__B1 _16451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24738__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13347__B1 _11626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21409__A1 _22501_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14255_ _14255_/A VGND VGND VPWR VPWR _14255_/Y sky130_fd_sc_hd__inv_2
X_17043_ _17128_/A _17043_/B _17040_/X _17042_/X VGND VGND VPWR VPWR _17044_/B sky130_fd_sc_hd__or4_4
XFILLER_7_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14206__A _14206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18901__A _18763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13206_ _13238_/A _13204_/X _13206_/C VGND VGND VPWR VPWR _13207_/C sky130_fd_sc_hd__and3_4
X_14186_ _24827_/Q _14169_/B _24826_/Q _14165_/B VGND VGND VPWR VPWR _14186_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23810__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24391__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22423__A _21569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13137_ _13137_/A _13137_/B VGND VGND VPWR VPWR _13138_/C sky130_fd_sc_hd__or2_4
X_18994_ _21940_/B _18991_/X _15545_/X _18991_/X VGND VGND VPWR VPWR _18994_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16421__A _16426_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24320__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13068_ _13300_/A _13068_/B VGND VGND VPWR VPWR _13068_/X sky130_fd_sc_hd__or2_4
X_17945_ _17817_/A _23143_/Q VGND VGND VPWR VPWR _17946_/C sky130_fd_sc_hd__or2_4
XANTENNA__21039__A _11516_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12019_ _11994_/Y _12019_/B VGND VGND VPWR VPWR _12019_/Y sky130_fd_sc_hd__nor2_4
X_17876_ _17708_/X _17875_/X _23929_/Q _17767_/X VGND VGND VPWR VPWR _23929_/D sky130_fd_sc_hd__o22a_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20878__A _21072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19615_ _21336_/B _19613_/X _19614_/X _19613_/X VGND VGND VPWR VPWR _23273_/D sky130_fd_sc_hd__a2bb2o_4
X_16827_ _16780_/Y _16784_/Y _16827_/C VGND VGND VPWR VPWR _16885_/A sky130_fd_sc_hd__or3_4
XANTENNA__15811__A2 _15439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19546_ _19533_/Y VGND VGND VPWR VPWR _19546_/X sky130_fd_sc_hd__buf_2
X_16758_ _16758_/A VGND VGND VPWR VPWR _16834_/D sky130_fd_sc_hd__inv_2
XFILLER_80_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15709_ _16216_/A VGND VGND VPWR VPWR _15709_/X sky130_fd_sc_hd__buf_2
X_19477_ _19477_/A VGND VGND VPWR VPWR _19477_/Y sky130_fd_sc_hd__inv_2
X_16689_ _15959_/Y _17498_/A _15959_/Y _17498_/A VGND VGND VPWR VPWR _16689_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_26_0_HCLK clkbuf_5_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_53_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18428_ _18517_/A VGND VGND VPWR VPWR _18518_/A sky130_fd_sc_hd__inv_2
XFILLER_94_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18359_ _24208_/Q _23831_/Q _16428_/Y _18358_/Y VGND VGND VPWR VPWR _18359_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22845__B1 _24528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21370_ _21392_/A _19457_/Y VGND VGND VPWR VPWR _21372_/B sky130_fd_sc_hd__or2_4
XANTENNA__20320__A1 _14255_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16524__B1 _16093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24479__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20321_ _20320_/X VGND VGND VPWR VPWR _20321_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24408__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23040_ _23040_/A _23039_/X VGND VGND VPWR VPWR _23040_/X sky130_fd_sc_hd__and2_4
X_20252_ _20252_/A _20194_/B _20252_/C _20252_/D VGND VGND VPWR VPWR _20252_/X sky130_fd_sc_hd__or4_4
XANTENNA__12010__B1 _11981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22333__A _21570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20183_ _20249_/A _20234_/B VGND VGND VPWR VPWR _20183_/X sky130_fd_sc_hd__and2_4
XANTENNA__24061__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23022__B1 _22858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24991_ _24841_/CLK _13347_/X HRESETn VGND VGND VPWR VPWR _24991_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22987__B _23020_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21891__B _22024_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23942_ _23972_/CLK _23942_/D HRESETn VGND VGND VPWR VPWR _20778_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20788__A _15653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23873_ _23767_/CLK _23873_/D HRESETn VGND VGND VPWR VPWR _23873_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22824_ _21030_/X _22823_/X _22646_/X _24420_/Q _22647_/X VGND VGND VPWR VPWR _22824_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_72_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22755_ _22754_/X VGND VGND VPWR VPWR _22755_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15015__B1 _15003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21706_ _21706_/A _21602_/X _21653_/X _21705_/X VGND VGND VPWR VPWR HRDATA[4] sky130_fd_sc_hd__or4_4
XFILLER_13_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22686_ _22686_/A _22686_/B _22686_/C VGND VGND VPWR VPWR _22686_/X sky130_fd_sc_hd__or3_4
XFILLER_9_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24425_ _24425_/CLK _24425_/D HRESETn VGND VGND VPWR VPWR _15830_/A sky130_fd_sc_hd__dfrtp_4
X_21637_ _21636_/X VGND VGND VPWR VPWR _21653_/B sky130_fd_sc_hd__inv_2
XFILLER_138_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19089__A _18678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16506__A _16499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15410__A _22024_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22227__B _22227_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12370_ _12415_/A _24490_/Q _12415_/A _24490_/Q VGND VGND VPWR VPWR _12376_/B sky130_fd_sc_hd__a2bb2o_4
X_24356_ _23469_/CLK _16036_/Y HRESETn VGND VGND VPWR VPWR _13473_/A sky130_fd_sc_hd__dfstp_4
X_21568_ _24549_/Q _21292_/X _21107_/X _21567_/X VGND VGND VPWR VPWR _21568_/X sky130_fd_sc_hd__a211o_4
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24831__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23307_ _23282_/CLK _23307_/D VGND VGND VPWR VPWR _19518_/A sky130_fd_sc_hd__dfxtp_4
X_20519_ _20511_/X _20518_/Y _15347_/A _20515_/X VGND VGND VPWR VPWR _23717_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20862__A2 _21093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24287_ _23353_/CLK _16227_/X HRESETn VGND VGND VPWR VPWR _14431_/A sky130_fd_sc_hd__dfrtp_4
X_21499_ _21235_/A _19000_/Y VGND VGND VPWR VPWR _21499_/X sky130_fd_sc_hd__or2_4
XFILLER_101_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24149__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_46_0_HCLK clkbuf_7_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_93_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_14040_ _14039_/Y _14037_/X _13398_/X _14027_/X VGND VGND VPWR VPWR _14040_/X sky130_fd_sc_hd__a2bb2o_4
X_23238_ _23246_/CLK _23238_/D VGND VGND VPWR VPWR _23238_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23169_ _25112_/CLK _19898_/X VGND VGND VPWR VPWR _23169_/Q sky130_fd_sc_hd__dfxtp_4
X_15991_ _15991_/A VGND VGND VPWR VPWR _15991_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12304__B2 _24478_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17730_ _17817_/A _23429_/Q VGND VGND VPWR VPWR _17731_/C sky130_fd_sc_hd__or2_4
X_14942_ _14941_/Y _24269_/Q _14941_/Y _24269_/Q VGND VGND VPWR VPWR _14943_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23784__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17661_ _13406_/B VGND VGND VPWR VPWR _17662_/B sky130_fd_sc_hd__inv_2
XFILLER_75_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14873_ _15059_/A _14873_/B _15058_/A _14873_/D VGND VGND VPWR VPWR _14878_/A sky130_fd_sc_hd__or4_4
X_19400_ _19399_/Y _19397_/X _19308_/X _19397_/X VGND VGND VPWR VPWR _23349_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23713__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16612_ _14801_/Y _16610_/X _16376_/X _16610_/X VGND VGND VPWR VPWR _16612_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13824_ _24907_/Q VGND VGND VPWR VPWR _13824_/X sky130_fd_sc_hd__buf_2
XFILLER_47_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12068__B1 _11981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17592_ _17486_/A _17590_/A VGND VGND VPWR VPWR _17593_/C sky130_fd_sc_hd__or2_4
X_19331_ _23373_/Q VGND VGND VPWR VPWR _19331_/Y sky130_fd_sc_hd__inv_2
X_16543_ _21729_/A _16542_/X _16376_/X _16542_/X VGND VGND VPWR VPWR _24163_/D sky130_fd_sc_hd__a2bb2o_4
X_13755_ _13773_/D _13737_/A VGND VGND VPWR VPWR _13769_/D sky130_fd_sc_hd__or2_4
XFILLER_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19940__B1 _15556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13105__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12706_ _12701_/A _12701_/B _12674_/X _12703_/B VGND VGND VPWR VPWR _12707_/A sky130_fd_sc_hd__a211o_4
X_19262_ _19258_/Y _19261_/X _19170_/X _19261_/X VGND VGND VPWR VPWR _19262_/X sky130_fd_sc_hd__a2bb2o_4
X_16474_ _16473_/Y _16395_/X _16219_/X _16395_/X VGND VGND VPWR VPWR _24190_/D sky130_fd_sc_hd__a2bb2o_4
X_13686_ _23688_/Q VGND VGND VPWR VPWR _13686_/X sky130_fd_sc_hd__buf_2
XFILLER_70_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22418__A _22163_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24919__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18213_ _18300_/A _18327_/A _18212_/Y _18213_/D VGND VGND VPWR VPWR _18213_/X sky130_fd_sc_hd__or4_4
X_15425_ _15424_/Y VGND VGND VPWR VPWR _20861_/B sky130_fd_sc_hd__buf_2
X_12637_ _12636_/X VGND VGND VPWR VPWR _12637_/X sky130_fd_sc_hd__buf_2
X_19193_ _23421_/Q VGND VGND VPWR VPWR _19193_/Y sky130_fd_sc_hd__inv_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15320__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18144_ _16125_/Y _23845_/Q _16125_/Y _23845_/Q VGND VGND VPWR VPWR _18145_/D sky130_fd_sc_hd__a2bb2o_4
X_12568_ _12568_/A VGND VGND VPWR VPWR _12647_/B sky130_fd_sc_hd__inv_2
X_15356_ _22624_/A _15353_/X _11566_/X _15353_/X VGND VGND VPWR VPWR _15356_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12240__B1 _12195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24572__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16135__B _16135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11519_ _11518_/Y VGND VGND VPWR VPWR _11599_/A sky130_fd_sc_hd__buf_2
X_14307_ _14306_/Y _14300_/X _14218_/X _14288_/A VGND VGND VPWR VPWR _24784_/D sky130_fd_sc_hd__a2bb2o_4
X_18075_ _18075_/A _11728_/X VGND VGND VPWR VPWR _18075_/X sky130_fd_sc_hd__or2_4
XFILLER_129_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12499_ _12509_/A _12499_/B _12499_/C VGND VGND VPWR VPWR _12499_/X sky130_fd_sc_hd__and3_4
X_15287_ _15284_/Y _15285_/X _15286_/X _15285_/X VGND VGND VPWR VPWR _15287_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20880__B _11725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24501__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17026_ _17026_/A _17026_/B VGND VGND VPWR VPWR _17045_/C sky130_fd_sc_hd__or2_4
X_14238_ _14234_/Y _14226_/X _14236_/X _14237_/X VGND VGND VPWR VPWR _24813_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14169_ _12048_/B _14169_/B VGND VGND VPWR VPWR _14170_/C sky130_fd_sc_hd__or2_4
XFILLER_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16151__A _24315_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_3_0_HCLK clkbuf_6_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__21992__A _22249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18977_ _13161_/B VGND VGND VPWR VPWR _18977_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15493__B1 _11573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17928_ _17928_/A _18754_/A VGND VGND VPWR VPWR _17929_/C sky130_fd_sc_hd__or2_4
XFILLER_38_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19462__A _15561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17234__A1 _17224_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17859_ _17955_/A _17851_/X _17859_/C VGND VGND VPWR VPWR _17859_/X sky130_fd_sc_hd__and3_4
X_20870_ _20826_/A VGND VGND VPWR VPWR _21638_/A sky130_fd_sc_hd__buf_2
XFILLER_121_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16993__B1 _16205_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19529_ _19529_/A VGND VGND VPWR VPWR _22094_/B sky130_fd_sc_hd__inv_2
XFILLER_74_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18806__A _13038_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22540_ _12592_/Y _22539_/X _12823_/Y _22029_/X VGND VGND VPWR VPWR _22540_/X sky130_fd_sc_hd__o22a_4
XFILLER_14_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22471_ _20748_/X _22468_/Y _21029_/X _22470_/X VGND VGND VPWR VPWR _22471_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22818__B1 _24527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16326__A _16339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22047__B _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24210_ _24262_/CLK _16424_/X HRESETn VGND VGND VPWR VPWR _24210_/Q sky130_fd_sc_hd__dfrtp_4
X_21422_ _16041_/X _21422_/B _21422_/C VGND VGND VPWR VPWR _21458_/A sky130_fd_sc_hd__and3_4
X_25190_ _23085_/CLK _25190_/D HRESETn VGND VGND VPWR VPWR _25190_/Q sky130_fd_sc_hd__dfrtp_4
X_24141_ _24145_/CLK _24141_/D HRESETn VGND VGND VPWR VPWR _14812_/A sky130_fd_sc_hd__dfrtp_4
X_21353_ _21130_/X _21353_/B _21353_/C VGND VGND VPWR VPWR _21353_/X sky130_fd_sc_hd__and3_4
XANTENNA__24242__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20304_ _14264_/Y _20296_/X _20287_/X _20303_/X VGND VGND VPWR VPWR _20305_/A sky130_fd_sc_hd__a211o_4
XFILLER_11_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24072_ _24088_/CLK _24072_/D HRESETn VGND VGND VPWR VPWR _16829_/A sky130_fd_sc_hd__dfrtp_4
X_21284_ _21019_/A VGND VGND VPWR VPWR _22610_/A sky130_fd_sc_hd__buf_2
X_23023_ _23023_/A _23023_/B _23022_/X VGND VGND VPWR VPWR _23030_/C sky130_fd_sc_hd__and3_4
X_20235_ _20188_/A _13891_/A _20193_/A _20235_/D VGND VGND VPWR VPWR _20235_/X sky130_fd_sc_hd__and4_4
XANTENNA__16061__A _16061_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20166_ _20162_/B VGND VGND VPWR VPWR _20249_/A sky130_fd_sc_hd__buf_2
XFILLER_39_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18017__A3 _11643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20097_ _20097_/A VGND VGND VPWR VPWR _20110_/A sky130_fd_sc_hd__inv_2
X_24974_ _24974_/CLK _24974_/D HRESETn VGND VGND VPWR VPWR _13396_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_58_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23925_ _23925_/CLK _23925_/D HRESETn VGND VGND VPWR VPWR _23925_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16579__A3 _15596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11870_ _11862_/Y _11648_/X _11867_/X _13053_/A _11869_/Y VGND VGND VPWR VPWR _25168_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25030__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12852__A2_N _24455_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23856_ _24879_/CLK _18309_/X HRESETn VGND VGND VPWR VPWR _18212_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15124__B _15123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22807_ _16061_/A _22549_/A _22581_/X VGND VGND VPWR VPWR _22807_/X sky130_fd_sc_hd__o21a_4
X_20999_ _21006_/A _18849_/Y VGND VGND VPWR VPWR _20999_/X sky130_fd_sc_hd__or2_4
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23787_ _24788_/CLK _20690_/X HRESETn VGND VGND VPWR VPWR _11884_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_38_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17620__A _17614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13540_ _13540_/A _13539_/X VGND VGND VPWR VPWR _13540_/X sky130_fd_sc_hd__or2_4
XFILLER_25_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22738_ _21569_/A _22738_/B _22738_/C VGND VGND VPWR VPWR _22743_/B sky130_fd_sc_hd__and3_4
XANTENNA__21142__A _21469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13471_ _13471_/A VGND VGND VPWR VPWR _13474_/A sky130_fd_sc_hd__inv_2
X_22669_ _22668_/X VGND VGND VPWR VPWR _22687_/B sky130_fd_sc_hd__inv_2
XFILLER_40_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12422_ _12434_/A _12422_/B _12421_/X VGND VGND VPWR VPWR _12422_/X sky130_fd_sc_hd__and3_4
X_15210_ _15108_/B _15213_/B VGND VGND VPWR VPWR _15210_/Y sky130_fd_sc_hd__nand2_4
XFILLER_138_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24408_ _24412_/CLK _24408_/D HRESETn VGND VGND VPWR VPWR _24408_/Q sky130_fd_sc_hd__dfrtp_4
X_16190_ _24300_/Q VGND VGND VPWR VPWR _16190_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19150__B2 _19146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12353_ _22565_/A VGND VGND VPWR VPWR _12353_/Y sky130_fd_sc_hd__inv_2
X_15141_ _14888_/Y _15139_/A VGND VGND VPWR VPWR _15141_/X sky130_fd_sc_hd__or2_4
XANTENNA__20835__A2 _20831_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24339_ _24222_/CLK _24339_/D HRESETn VGND VGND VPWR VPWR _24339_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15072_ _14743_/X _15075_/B _14984_/X VGND VGND VPWR VPWR _15072_/Y sky130_fd_sc_hd__a21oi_4
X_12284_ _12165_/X VGND VGND VPWR VPWR _12300_/C sky130_fd_sc_hd__buf_2
XANTENNA__22037__B2 _21357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14023_ _13711_/X _23690_/Q VGND VGND VPWR VPWR _14023_/X sky130_fd_sc_hd__or2_4
X_18900_ _18899_/Y VGND VGND VPWR VPWR _18900_/X sky130_fd_sc_hd__buf_2
XFILLER_107_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17067__A _17067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19880_ _19880_/A VGND VGND VPWR VPWR _21008_/B sky130_fd_sc_hd__inv_2
XFILLER_134_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21796__B1 _21582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18831_ _14548_/X _14549_/X _14539_/Y _19862_/B VGND VGND VPWR VPWR _18832_/A sky130_fd_sc_hd__or4_4
XANTENNA__23965__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_133_0_HCLK clkbuf_7_66_0_HCLK/X VGND VGND VPWR VPWR _23586_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__25189__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_196_0_HCLK clkbuf_7_98_0_HCLK/X VGND VGND VPWR VPWR _23702_/CLK sky130_fd_sc_hd__clkbuf_1
X_18762_ _18776_/A VGND VGND VPWR VPWR _18762_/X sky130_fd_sc_hd__buf_2
X_15974_ _15972_/Y _15973_/X _11598_/X _15973_/X VGND VGND VPWR VPWR _24371_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25118__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21548__B1 _21546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22420__B _22147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17713_ _17729_/A VGND VGND VPWR VPWR _17853_/A sky130_fd_sc_hd__buf_2
X_14925_ _14925_/A VGND VGND VPWR VPWR _15110_/B sky130_fd_sc_hd__inv_2
X_18693_ _18689_/Y _18692_/X _17199_/X _18692_/X VGND VGND VPWR VPWR _23598_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17644_ _17644_/A VGND VGND VPWR VPWR _21144_/A sky130_fd_sc_hd__buf_2
XFILLER_63_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14856_ _15064_/A _16601_/A _24686_/Q _14835_/Y VGND VGND VPWR VPWR _14856_/X sky130_fd_sc_hd__a2bb2o_4
X_13807_ _13806_/X VGND VGND VPWR VPWR _13811_/B sky130_fd_sc_hd__inv_2
X_17575_ _17497_/B _17548_/X _17520_/X _17572_/B VGND VGND VPWR VPWR _17575_/X sky130_fd_sc_hd__a211o_4
X_14787_ _24712_/Q VGND VGND VPWR VPWR _14977_/C sky130_fd_sc_hd__inv_2
X_11999_ _11999_/A VGND VGND VPWR VPWR _11999_/Y sky130_fd_sc_hd__inv_2
X_19314_ _13178_/B VGND VGND VPWR VPWR _19314_/Y sky130_fd_sc_hd__inv_2
X_16526_ _22343_/A _16523_/X _16096_/X _16523_/X VGND VGND VPWR VPWR _16526_/X sky130_fd_sc_hd__a2bb2o_4
X_13738_ _13722_/X _13745_/B _13745_/A _13725_/Y VGND VGND VPWR VPWR _13738_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22148__A _22148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24753__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19245_ _21826_/B _19239_/X _11844_/X _19244_/X VGND VGND VPWR VPWR _23404_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21052__A _21051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16457_ _16457_/A VGND VGND VPWR VPWR _16457_/Y sky130_fd_sc_hd__inv_2
X_13669_ _13428_/Y _13667_/X _13668_/X _13667_/X VGND VGND VPWR VPWR _24930_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15408_ _15407_/Y VGND VGND VPWR VPWR _21113_/B sky130_fd_sc_hd__buf_2
X_19176_ _19174_/Y _19169_/X _19152_/X _19175_/X VGND VGND VPWR VPWR _19176_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21987__A _21292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16388_ _16387_/Y _16308_/A _16219_/X _16308_/A VGND VGND VPWR VPWR _24222_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18127_ _18127_/A VGND VGND VPWR VPWR _18127_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13961__B1 _24805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15339_ _15339_/A VGND VGND VPWR VPWR _22810_/A sky130_fd_sc_hd__inv_2
XFILLER_129_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21577__A2_N _21576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18058_ _18023_/X _17640_/Y _18023_/X _17640_/Y VGND VGND VPWR VPWR _18058_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14505__A2 _14480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12516__A1 _12345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20039__B1 _19714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17009_ _16151_/Y _24053_/Q _24309_/Q _17097_/A VGND VGND VPWR VPWR _17012_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_92_0_HCLK clkbuf_6_46_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_92_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20020_ _20014_/Y VGND VGND VPWR VPWR _20020_/X sky130_fd_sc_hd__buf_2
XFILLER_8_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14269__B2 _14268_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12315__A1_N _12474_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23635__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18404__B1 _16464_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21971_ _20814_/X VGND VGND VPWR VPWR _22702_/A sky130_fd_sc_hd__buf_2
XFILLER_132_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22751__A2 _21553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20922_ _20413_/A _11940_/Y _20740_/B _21638_/A VGND VGND VPWR VPWR _20922_/X sky130_fd_sc_hd__o22a_4
X_23710_ _23744_/CLK _23710_/D HRESETn VGND VGND VPWR VPWR _13509_/A sky130_fd_sc_hd__dfrtp_4
X_24690_ _24264_/CLK _15075_/X HRESETn VGND VGND VPWR VPWR _24690_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20762__B2 _15642_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20853_ _11503_/A VGND VGND VPWR VPWR _21432_/A sky130_fd_sc_hd__buf_2
XPHY_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23641_ _23641_/CLK _20328_/Y HRESETn VGND VGND VPWR VPWR _18619_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23572_ _23560_/CLK _18770_/X VGND VGND VPWR VPWR _18768_/A sky130_fd_sc_hd__dfxtp_4
X_20784_ _20783_/X VGND VGND VPWR VPWR _22501_/A sky130_fd_sc_hd__buf_2
XANTENNA__21711__B1 _24400_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24494__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22523_ _22522_/X VGND VGND VPWR VPWR _22523_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16056__A _16056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24423__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22454_ _22219_/A _22451_/X _20750_/X _22453_/X VGND VGND VPWR VPWR _22455_/A sky130_fd_sc_hd__o22a_4
XFILLER_10_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21405_ _21404_/X VGND VGND VPWR VPWR _21405_/Y sky130_fd_sc_hd__inv_2
X_25173_ _23246_/CLK _25173_/D HRESETn VGND VGND VPWR VPWR _11842_/A sky130_fd_sc_hd__dfrtp_4
X_22385_ _22385_/A _20787_/B VGND VGND VPWR VPWR _22385_/X sky130_fd_sc_hd__or2_4
XFILLER_108_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24124_ _24094_/CLK _16623_/X HRESETn VGND VGND VPWR VPWR _24124_/Q sky130_fd_sc_hd__dfrtp_4
X_21336_ _21336_/A _21336_/B VGND VGND VPWR VPWR _21337_/C sky130_fd_sc_hd__or2_4
XANTENNA__22019__B2 _21408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24055_ _24055_/CLK _17066_/Y HRESETn VGND VGND VPWR VPWR _24055_/Q sky130_fd_sc_hd__dfrtp_4
X_21267_ _21042_/X _21266_/X _21046_/X _25192_/Q _21047_/X VGND VGND VPWR VPWR _21268_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_137_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14304__A _16216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16222__C _16222_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23006_ _23026_/B _23005_/X _22459_/X _24533_/Q _22460_/X VGND VGND VPWR VPWR _23006_/X
+ sky130_fd_sc_hd__a32o_4
X_20218_ _20245_/A _20210_/X _20217_/Y VGND VGND VPWR VPWR _20241_/A sky130_fd_sc_hd__o21a_4
XFILLER_46_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21198_ _20994_/A VGND VGND VPWR VPWR _21234_/A sky130_fd_sc_hd__buf_2
XFILLER_103_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_206_0_HCLK clkbuf_8_207_0_HCLK/A VGND VGND VPWR VPWR _23706_/CLK sky130_fd_sc_hd__clkbuf_1
X_20149_ _20147_/Y _20148_/X _19808_/X _20148_/X VGND VGND VPWR VPWR _23071_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17615__A _17615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25211__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21137__A _21469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12971_ _12933_/C _12878_/C VGND VGND VPWR VPWR _12972_/B sky130_fd_sc_hd__or2_4
X_24957_ _24957_/CLK _13584_/X HRESETn VGND VGND VPWR VPWR _11673_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14710_ _24708_/Q VGND VGND VPWR VPWR _14880_/A sky130_fd_sc_hd__inv_2
X_11922_ _21897_/A _11919_/X _11923_/A _11919_/X VGND VGND VPWR VPWR _25163_/D sky130_fd_sc_hd__a2bb2o_4
X_23908_ _23908_/CLK _23908_/D HRESETn VGND VGND VPWR VPWR _23908_/Q sky130_fd_sc_hd__dfrtp_4
X_15690_ _15684_/X _15689_/X _16093_/A _24480_/Q _15685_/X VGND VGND VPWR VPWR _24480_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24800__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24888_ _23774_/CLK _13979_/X HRESETn VGND VGND VPWR VPWR _24888_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14641_ _14643_/A _14638_/X _14639_/Y _14640_/X VGND VGND VPWR VPWR _14641_/X sky130_fd_sc_hd__o22a_4
XFILLER_122_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24863__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11853_ _19610_/A VGND VGND VPWR VPWR _11853_/X sky130_fd_sc_hd__buf_2
X_23839_ _23826_/CLK _23839_/D HRESETn VGND VGND VPWR VPWR _23839_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17360_ _17306_/Y _17362_/B _17359_/Y VGND VGND VPWR VPWR _17360_/X sky130_fd_sc_hd__o21a_4
XFILLER_92_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11784_ _17448_/B _11784_/B _11783_/X VGND VGND VPWR VPWR _11803_/C sky130_fd_sc_hd__and3_4
X_14572_ _14571_/X VGND VGND VPWR VPWR _14573_/A sky130_fd_sc_hd__buf_2
XFILLER_13_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12443__B1 _12416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16311_ _16310_/Y _16308_/X _16141_/X _16308_/X VGND VGND VPWR VPWR _24252_/D sky130_fd_sc_hd__a2bb2o_4
X_13523_ _20635_/A _20635_/B _20635_/C _23746_/Q VGND VGND VPWR VPWR _13524_/D sky130_fd_sc_hd__or4_4
X_17291_ _11628_/Y _17318_/A _25191_/Q _17323_/C VGND VGND VPWR VPWR _17291_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24164__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19030_ _20998_/B _19025_/X _18662_/X _19012_/Y VGND VGND VPWR VPWR _23479_/D sky130_fd_sc_hd__a2bb2o_4
X_16242_ _16247_/A VGND VGND VPWR VPWR _16242_/X sky130_fd_sc_hd__buf_2
X_13454_ _13454_/A _13427_/X _13440_/X _13453_/X VGND VGND VPWR VPWR _13454_/X sky130_fd_sc_hd__or4_4
XFILLER_103_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12405_ _12388_/Y _12534_/A _12536_/A _12405_/D VGND VGND VPWR VPWR _12409_/C sky130_fd_sc_hd__or4_4
XANTENNA__21600__A _21585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13385_ _11916_/X VGND VGND VPWR VPWR _20686_/B sky130_fd_sc_hd__inv_2
X_16173_ _16172_/Y _16170_/X _15775_/X _16170_/X VGND VGND VPWR VPWR _24307_/D sky130_fd_sc_hd__a2bb2o_4
X_15124_ _15117_/X _15123_/X VGND VGND VPWR VPWR _15125_/B sky130_fd_sc_hd__or2_4
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12336_ _25077_/Q _24474_/Q _12407_/B _12335_/Y VGND VGND VPWR VPWR _12336_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15696__B1 _13658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_16_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_16_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_12267_ _12180_/A _12267_/B VGND VGND VPWR VPWR _12283_/B sky130_fd_sc_hd__or2_4
X_15055_ _15019_/B _15049_/X _15027_/X _15051_/Y VGND VGND VPWR VPWR _15055_/X sky130_fd_sc_hd__a211o_4
X_19932_ _19926_/Y VGND VGND VPWR VPWR _19932_/X sky130_fd_sc_hd__buf_2
X_14006_ _14004_/Y _13937_/X _13963_/X _14005_/Y VGND VGND VPWR VPWR _14007_/A sky130_fd_sc_hd__o22a_4
X_19863_ _19863_/A VGND VGND VPWR VPWR _19876_/A sky130_fd_sc_hd__inv_2
XANTENNA__18634__B1 _16556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12198_ _12170_/B _12186_/B _12192_/A VGND VGND VPWR VPWR _12198_/X sky130_fd_sc_hd__or3_4
XFILLER_68_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18814_ _18809_/A VGND VGND VPWR VPWR _18814_/X sky130_fd_sc_hd__buf_2
XANTENNA__17525__A _16693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19794_ _19792_/Y _19793_/X _19459_/X _19793_/X VGND VGND VPWR VPWR _19794_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18745_ _18752_/A VGND VGND VPWR VPWR _18745_/X sky130_fd_sc_hd__buf_2
XFILLER_49_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15957_ _15957_/A VGND VGND VPWR VPWR _15957_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13675__A1_N _13441_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22733__A2 _22281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11573__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14908_ _24669_/Q _24274_/Q _15105_/A _14907_/Y VGND VGND VPWR VPWR _14918_/A sky130_fd_sc_hd__o22a_4
XANTENNA__15045__A _15045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18676_ _18675_/Y _18673_/X _16546_/X _18673_/X VGND VGND VPWR VPWR _23603_/D sky130_fd_sc_hd__a2bb2o_4
X_15888_ _15887_/Y _15885_/X _15513_/X _15885_/X VGND VGND VPWR VPWR _15888_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24934__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17627_ _17626_/X VGND VGND VPWR VPWR _17648_/B sky130_fd_sc_hd__inv_2
X_14839_ _24692_/Q VGND VGND VPWR VPWR _14839_/Y sky130_fd_sc_hd__inv_2
X_17558_ _16697_/Y _17558_/B _17498_/Y _17550_/B VGND VGND VPWR VPWR _17564_/B sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_5_26_0_HCLK_A clkbuf_5_27_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18075__B _11728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16509_ _16508_/Y _16506_/X _16261_/X _16506_/X VGND VGND VPWR VPWR _16509_/X sky130_fd_sc_hd__a2bb2o_4
X_17489_ _17487_/Y _17615_/A _17489_/C _17488_/Y VGND VGND VPWR VPWR _17489_/X sky130_fd_sc_hd__or4_4
XFILLER_108_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19228_ _19225_/Y _19226_/X _19227_/X _19226_/X VGND VGND VPWR VPWR _19228_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22606__A _22178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21510__A _21394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19159_ _17884_/B VGND VGND VPWR VPWR _19159_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23887__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22170_ _21020_/B VGND VGND VPWR VPWR _22170_/X sky130_fd_sc_hd__buf_2
XANTENNA__15687__B1 _24482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21121_ SSn_S3 _11952_/X _21179_/A VGND VGND VPWR VPWR _21121_/X sky130_fd_sc_hd__o21a_4
XANTENNA__23816__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21052_ _21051_/X VGND VGND VPWR VPWR _22245_/A sky130_fd_sc_hd__buf_2
XANTENNA__22421__A1 _24516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20003_ _19990_/Y VGND VGND VPWR VPWR _20003_/X sky130_fd_sc_hd__buf_2
XFILLER_87_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22060__B _19486_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24811_ _24811_/CLK _14242_/X HRESETn VGND VGND VPWR VPWR _24811_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__22185__B1 _24554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_36_0_HCLK clkbuf_8_37_0_HCLK/A VGND VGND VPWR VPWR _23249_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__19050__B1 _18959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24742_ _25106_/CLK _14545_/Y HRESETn VGND VGND VPWR VPWR _24742_/Q sky130_fd_sc_hd__dfrtp_4
X_21954_ _21378_/A _19783_/Y VGND VGND VPWR VPWR _21955_/C sky130_fd_sc_hd__or2_4
Xclkbuf_8_99_0_HCLK clkbuf_8_99_0_HCLK/A VGND VGND VPWR VPWR _24064_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24675__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20905_ _21716_/B _20904_/X _23040_/A _22859_/A VGND VGND VPWR VPWR _20905_/X sky130_fd_sc_hd__o22a_4
XPHY_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21885_ _25144_/Q _21881_/Y _21883_/X _21884_/Y VGND VGND VPWR VPWR _21885_/X sky130_fd_sc_hd__a211o_4
XFILLER_55_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24673_ _24676_/CLK _24673_/D HRESETn VGND VGND VPWR VPWR _24673_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24604__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15105__D _14941_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _20820_/X _20822_/Y _20835_/X VGND VGND VPWR VPWR _20836_/X sky130_fd_sc_hd__and3_4
XPHY_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23624_ _23624_/CLK _23624_/D HRESETn VGND VGND VPWR VPWR _23624_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20767_ _20931_/A VGND VGND VPWR VPWR _22445_/B sky130_fd_sc_hd__buf_2
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23555_ _23133_/CLK _18818_/X VGND VGND VPWR VPWR _13156_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_50_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17320__D _17415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22506_ _24340_/Q _22350_/X _22351_/X VGND VGND VPWR VPWR _22506_/X sky130_fd_sc_hd__o21a_4
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15914__A1 _11535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23486_ _23486_/CLK _23486_/D VGND VGND VPWR VPWR _23486_/Q sky130_fd_sc_hd__dfxtp_4
X_20698_ _20698_/A _20697_/B VGND VGND VPWR VPWR _20698_/X sky130_fd_sc_hd__and2_4
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22437_ _11583_/A _22435_/X _20744_/X _22436_/X VGND VGND VPWR VPWR _22437_/X sky130_fd_sc_hd__a211o_4
XFILLER_104_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13170_ _13301_/A _13170_/B VGND VGND VPWR VPWR _13171_/C sky130_fd_sc_hd__or2_4
X_22368_ _21978_/X _22367_/X VGND VGND VPWR VPWR _22368_/X sky130_fd_sc_hd__and2_4
XANTENNA__18864__B1 _18795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25156_ _24088_/CLK _11958_/X HRESETn VGND VGND VPWR VPWR _25156_/Q sky130_fd_sc_hd__dfrtp_4
X_12121_ _24562_/Q VGND VGND VPWR VPWR _12121_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15678__B1 _15350_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21319_ _17615_/A _11514_/X _12818_/Y _15576_/X VGND VGND VPWR VPWR _21319_/X sky130_fd_sc_hd__o22a_4
X_24107_ _24112_/CLK _16654_/X HRESETn VGND VGND VPWR VPWR _24107_/Q sky130_fd_sc_hd__dfrtp_4
X_25087_ _25091_/CLK _12483_/X HRESETn VGND VGND VPWR VPWR _22564_/A sky130_fd_sc_hd__dfrtp_4
X_22299_ _22299_/A _22298_/X VGND VGND VPWR VPWR _22299_/X sky130_fd_sc_hd__and2_4
XANTENNA__17048__C _17067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13153__A1 _11711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12052_ _25137_/Q _20695_/B _12051_/X VGND VGND VPWR VPWR _12052_/X sky130_fd_sc_hd__a21o_4
XFILLER_78_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24038_ _24037_/CLK _24038_/D HRESETn VGND VGND VPWR VPWR _24038_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22412__B2 _22285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20423__B1 _20419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16860_ _16859_/X VGND VGND VPWR VPWR _24087_/D sky130_fd_sc_hd__inv_2
XFILLER_137_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15811_ _15720_/X _15439_/X _15712_/A _13456_/A VGND VGND VPWR VPWR _15811_/X sky130_fd_sc_hd__a211o_4
X_16791_ _16785_/X _16791_/B _16789_/X _16790_/X VGND VGND VPWR VPWR _16791_/X sky130_fd_sc_hd__or4_4
XFILLER_92_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12489__A _12489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18530_ _18540_/A _18530_/B _18530_/C VGND VGND VPWR VPWR _23824_/D sky130_fd_sc_hd__and3_4
XANTENNA__15850__B1 _11555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15742_ _15421_/X _15740_/X _15735_/X _24461_/Q _15741_/X VGND VGND VPWR VPWR _15742_/X
+ sky130_fd_sc_hd__a32o_4
X_12954_ _12953_/X VGND VGND VPWR VPWR _25021_/D sky130_fd_sc_hd__inv_2
XFILLER_133_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11905_ _11905_/A _11884_/X VGND VGND VPWR VPWR _11905_/X sky130_fd_sc_hd__and2_4
X_18461_ _23840_/Q _18466_/B VGND VGND VPWR VPWR _18461_/X sky130_fd_sc_hd__or2_4
X_15673_ _15658_/X _15672_/X _15596_/X _24492_/Q _15661_/X VGND VGND VPWR VPWR _15673_/X
+ sky130_fd_sc_hd__a32o_4
X_12885_ _12788_/Y _12884_/X VGND VGND VPWR VPWR _12885_/X sky130_fd_sc_hd__or2_4
XANTENNA__24345__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_7_0_HCLK clkbuf_5_6_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15602__B1 _11558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17412_ _17317_/C _17412_/B VGND VGND VPWR VPWR _17413_/B sky130_fd_sc_hd__or2_4
XFILLER_45_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14624_ _14633_/A _14610_/B _24719_/Q VGND VGND VPWR VPWR _14625_/B sky130_fd_sc_hd__or3_4
X_11836_ _11834_/Y _11831_/X _11835_/X _11831_/X VGND VGND VPWR VPWR _25175_/D sky130_fd_sc_hd__a2bb2o_4
X_18392_ _16436_/Y _18509_/A _16436_/Y _18509_/A VGND VGND VPWR VPWR _18392_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21314__B _21448_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17260_/Y _17340_/X VGND VGND VPWR VPWR _17343_/X sky130_fd_sc_hd__or2_4
X_14555_ _21257_/A _16035_/B _13462_/A VGND VGND VPWR VPWR _14555_/X sky130_fd_sc_hd__o21a_4
X_11767_ _11766_/Y VGND VGND VPWR VPWR _11767_/X sky130_fd_sc_hd__buf_2
XPHY_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _13506_/A _13506_/B _13506_/C _13506_/D VGND VGND VPWR VPWR _13506_/X sky130_fd_sc_hd__or4_4
XFILLER_18_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17274_ _25191_/Q _17323_/C _25195_/Q _17273_/Y VGND VGND VPWR VPWR _17274_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14486_ _14485_/Y VGND VGND VPWR VPWR _14486_/X sky130_fd_sc_hd__buf_2
X_11698_ _11645_/X _11697_/Y _11698_/C _11698_/D VGND VGND VPWR VPWR _11698_/X sky130_fd_sc_hd__and4_4
X_19013_ _19012_/Y VGND VGND VPWR VPWR _19013_/X sky130_fd_sc_hd__buf_2
X_16225_ _16224_/X VGND VGND VPWR VPWR _16225_/Y sky130_fd_sc_hd__inv_2
X_13437_ _24933_/Q VGND VGND VPWR VPWR _13437_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23980__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16156_ _16155_/Y _16152_/X _15479_/X _16152_/X VGND VGND VPWR VPWR _16156_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21454__A2 _15456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18855__B1 _18764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13368_ _13368_/A VGND VGND VPWR VPWR _21884_/A sky130_fd_sc_hd__inv_2
XFILLER_5_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15107_ _15104_/Y _15161_/A _15107_/C VGND VGND VPWR VPWR _15115_/A sky130_fd_sc_hd__or3_4
XFILLER_127_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12319_ _24488_/Q VGND VGND VPWR VPWR _12319_/Y sky130_fd_sc_hd__inv_2
X_16087_ _16087_/A VGND VGND VPWR VPWR _16087_/X sky130_fd_sc_hd__buf_2
XANTENNA__25133__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13299_ _13299_/A _13297_/X _13298_/X VGND VGND VPWR VPWR _13303_/B sky130_fd_sc_hd__and3_4
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15038_ _24699_/Q _15038_/B VGND VGND VPWR VPWR _15039_/C sky130_fd_sc_hd__or2_4
X_19915_ _19915_/A VGND VGND VPWR VPWR _21518_/B sky130_fd_sc_hd__inv_2
XFILLER_25_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22954__A2 _22281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14892__B2 _24280_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17285__A1_N _11623_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19846_ _23188_/Q VGND VGND VPWR VPWR _21774_/B sky130_fd_sc_hd__inv_2
XANTENNA__19280__B1 _19232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16094__B1 _16093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16989_ _21293_/A _21291_/A _16213_/Y _17161_/A VGND VGND VPWR VPWR _16989_/X sky130_fd_sc_hd__o22a_4
X_19777_ _19776_/Y _19772_/X _19755_/X _19759_/Y VGND VGND VPWR VPWR _23215_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_252_0_HCLK clkbuf_8_253_0_HCLK/A VGND VGND VPWR VPWR _24674_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18728_ _17920_/B VGND VGND VPWR VPWR _18728_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21505__A _21374_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18659_ _23608_/Q VGND VGND VPWR VPWR _18659_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24086__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15503__A _11532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21670_ _21675_/A _21668_/X _21669_/X VGND VGND VPWR VPWR _21670_/X sky130_fd_sc_hd__and3_4
XFILLER_40_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24015__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20621_ _20647_/A VGND VGND VPWR VPWR _20621_/X sky130_fd_sc_hd__buf_2
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17346__B1 _17345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23340_ _23350_/CLK _23340_/D VGND VGND VPWR VPWR _23340_/Q sky130_fd_sc_hd__dfxtp_4
X_20552_ _20601_/A VGND VGND VPWR VPWR _20552_/X sky130_fd_sc_hd__buf_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22336__A _24105_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21240__A _21393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23271_ _23356_/CLK _23271_/D VGND VGND VPWR VPWR _19619_/A sky130_fd_sc_hd__dfxtp_4
X_20483_ _20461_/X _20482_/X _24598_/Q _20466_/X VGND VGND VPWR VPWR _20483_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16334__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22222_ _22500_/A _22213_/X _22221_/X VGND VGND VPWR VPWR _22222_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_118_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17649__A1 _21144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25010_ _25012_/CLK _25010_/D HRESETn VGND VGND VPWR VPWR _25010_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22642__A1 _22369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23650__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22153_ _16366_/Y _22153_/B VGND VGND VPWR VPWR _22155_/B sky130_fd_sc_hd__or2_4
XFILLER_106_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19249__A2_N _19244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21104_ _21104_/A _21565_/A VGND VGND VPWR VPWR _21104_/X sky130_fd_sc_hd__and2_4
XFILLER_86_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22084_ _22084_/A _22084_/B VGND VGND VPWR VPWR _22084_/X sky130_fd_sc_hd__or2_4
XFILLER_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15675__A3 _15600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_62_0_HCLK clkbuf_6_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_62_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21035_ _21034_/Y VGND VGND VPWR VPWR _22646_/A sky130_fd_sc_hd__buf_2
XFILLER_114_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17165__A _17086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16085__B1 _11576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24856__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22986_ _22334_/A _22983_/X _22986_/C VGND VGND VPWR VPWR _22997_/B sky130_fd_sc_hd__and3_4
XFILLER_16_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24725_ _23661_/CLK _14656_/X HRESETn VGND VGND VPWR VPWR _24725_/Q sky130_fd_sc_hd__dfrtp_4
X_21937_ _21172_/X _21933_/X _21936_/X VGND VGND VPWR VPWR _21937_/X sky130_fd_sc_hd__or3_4
XFILLER_28_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11941__A _11940_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12670_ _12672_/B VGND VGND VPWR VPWR _12671_/B sky130_fd_sc_hd__inv_2
XFILLER_128_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24656_ _24662_/CLK _24656_/D HRESETn VGND VGND VPWR VPWR _14969_/A sky130_fd_sc_hd__dfrtp_4
X_21868_ _16539_/Y _21868_/B VGND VGND VPWR VPWR _21868_/X sky130_fd_sc_hd__and2_4
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18129__A2 _18112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11599_/A VGND VGND VPWR VPWR _11621_/X sky130_fd_sc_hd__buf_2
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23607_ _25050_/CLK _18663_/X VGND VGND VPWR VPWR _18661_/A sky130_fd_sc_hd__dfxtp_4
X_20819_ _20818_/X VGND VGND VPWR VPWR _20819_/X sky130_fd_sc_hd__buf_2
XFILLER_93_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21799_ _21799_/A _21181_/A VGND VGND VPWR VPWR _21799_/X sky130_fd_sc_hd__and2_4
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24587_ _24587_/CLK _24587_/D HRESETn VGND VGND VPWR VPWR _24587_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ _21443_/A _14325_/A _24774_/Q _14319_/X VGND VGND VPWR VPWR _14340_/X sky130_fd_sc_hd__o22a_4
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ HWDATA[24] VGND VGND VPWR VPWR _11552_/X sky130_fd_sc_hd__buf_2
XANTENNA__22881__A1 _16056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23538_ _23133_/CLK _18864_/X VGND VGND VPWR VPWR _18863_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16447__A1_N _16445_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22246__A _16193_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24631__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23738__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14271_ _14270_/Y _14268_/X _14232_/X _14268_/X VGND VGND VPWR VPWR _24798_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16560__A1 _15430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23469_ _23469_/CLK _19062_/X VGND VGND VPWR VPWR _17719_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_7_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16010_ _15439_/X _14435_/D _16005_/X _16008_/X _16009_/X VGND VGND VPWR VPWR _16011_/A
+ sky130_fd_sc_hd__o32a_4
X_13222_ _13222_/A _13218_/X _13222_/C VGND VGND VPWR VPWR _13222_/X sky130_fd_sc_hd__or3_4
X_25208_ _25012_/CLK _25208_/D HRESETn VGND VGND VPWR VPWR _11568_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21436__A2 _24258_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13153_ _11711_/X _13134_/X _13152_/X _25002_/Q _13114_/X VGND VGND VPWR VPWR _13153_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_83_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25139_ _24840_/CLK _25139_/D HRESETn VGND VGND VPWR VPWR _25139_/Q sky130_fd_sc_hd__dfrtp_4
X_12104_ _24552_/Q VGND VGND VPWR VPWR _12104_/Y sky130_fd_sc_hd__inv_2
X_13084_ _13169_/A VGND VGND VPWR VPWR _13085_/A sky130_fd_sc_hd__buf_2
X_17961_ _17961_/A _17959_/X _17960_/X VGND VGND VPWR VPWR _17961_/X sky130_fd_sc_hd__and3_4
XFILLER_97_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14699__A _24099_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22397__B1 _24040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12035_ _23798_/Q _12016_/X VGND VGND VPWR VPWR _12035_/X sky130_fd_sc_hd__and2_4
X_16912_ _16879_/A _16838_/X VGND VGND VPWR VPWR _16912_/X sky130_fd_sc_hd__or2_4
X_19700_ _23241_/Q VGND VGND VPWR VPWR _19700_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19262__B1 _19170_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17892_ _17924_/A _23569_/Q VGND VGND VPWR VPWR _17894_/B sky130_fd_sc_hd__or2_4
XFILLER_61_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21309__B _21097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24597__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16843_ _16879_/A _16774_/Y _16853_/A _16852_/B VGND VGND VPWR VPWR _16843_/X sky130_fd_sc_hd__or4_4
X_19631_ _19631_/A VGND VGND VPWR VPWR _21615_/B sky130_fd_sc_hd__inv_2
XFILLER_19_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24526__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19562_ _23291_/Q VGND VGND VPWR VPWR _21624_/B sky130_fd_sc_hd__inv_2
X_16774_ _16774_/A VGND VGND VPWR VPWR _16774_/Y sky130_fd_sc_hd__inv_2
X_13986_ _13926_/C _13941_/B _13926_/C _13941_/B VGND VGND VPWR VPWR _13986_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18513_ _18513_/A VGND VGND VPWR VPWR _18513_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15725_ _15717_/B _15722_/C VGND VGND VPWR VPWR _15726_/A sky130_fd_sc_hd__or2_4
X_12937_ _12937_/A VGND VGND VPWR VPWR _12937_/Y sky130_fd_sc_hd__inv_2
X_19493_ _19493_/A VGND VGND VPWR VPWR _19493_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12947__A _12947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_82_0_HCLK clkbuf_8_83_0_HCLK/A VGND VGND VPWR VPWR _24884_/CLK sky130_fd_sc_hd__clkbuf_1
X_18444_ _18463_/A _18444_/B _18443_/Y VGND VGND VPWR VPWR _23844_/D sky130_fd_sc_hd__and3_4
X_15656_ _22147_/A VGND VGND VPWR VPWR _15692_/A sky130_fd_sc_hd__buf_2
XANTENNA__21044__B _21043_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12868_ _12867_/X VGND VGND VPWR VPWR _12921_/A sky130_fd_sc_hd__buf_2
X_14607_ scl_oen_o_S5 _20729_/B _23665_/Q VGND VGND VPWR VPWR _14618_/B sky130_fd_sc_hd__and3_4
X_11819_ _11777_/A _11817_/X _11818_/Y VGND VGND VPWR VPWR _25179_/D sky130_fd_sc_hd__o21a_4
X_18375_ _23815_/Q VGND VGND VPWR VPWR _18552_/A sky130_fd_sc_hd__inv_2
X_15587_ _15574_/X _15582_/X _15468_/X _24532_/Q _15585_/X VGND VGND VPWR VPWR _15587_/X
+ sky130_fd_sc_hd__a32o_4
X_12799_ _22160_/A VGND VGND VPWR VPWR _12984_/A sky130_fd_sc_hd__inv_2
XPHY_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20883__B _15426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17326_ _17348_/D _17348_/B VGND VGND VPWR VPWR _17327_/D sky130_fd_sc_hd__or2_4
X_14538_ _14524_/B _14521_/X _14536_/X VGND VGND VPWR VPWR _24743_/D sky130_fd_sc_hd__o21a_4
XFILLER_30_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22872__A1 _13337_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_2_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_2_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__16000__B1 _15709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17257_ _17257_/A VGND VGND VPWR VPWR _17317_/C sky130_fd_sc_hd__inv_2
X_14469_ _24746_/Q VGND VGND VPWR VPWR _14469_/X sky130_fd_sc_hd__buf_2
X_16208_ _16137_/A VGND VGND VPWR VPWR _16208_/X sky130_fd_sc_hd__buf_2
XFILLER_127_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21995__A _22992_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17188_ _17187_/X VGND VGND VPWR VPWR _17188_/X sky130_fd_sc_hd__buf_2
X_16139_ _16133_/Y _16138_/X _15828_/X _16138_/X VGND VGND VPWR VPWR _24320_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18056__A1 _17446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20938__A1 _23025_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16067__B1 _11555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19829_ _21525_/B _19822_/X _19828_/X _19822_/X VGND VGND VPWR VPWR _19829_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24267__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22840_ _22840_/A VGND VGND VPWR VPWR _22840_/X sky130_fd_sc_hd__buf_2
XFILLER_77_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21235__A _21235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19556__B2 _19555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22771_ _17481_/A _22654_/X _22608_/X VGND VGND VPWR VPWR _22773_/C sky130_fd_sc_hd__a21o_4
XFILLER_52_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24510_ _25034_/CLK _15625_/X HRESETn VGND VGND VPWR VPWR _24510_/Q sky130_fd_sc_hd__dfrtp_4
X_21722_ _21715_/X _21717_/X _22547_/A _21721_/X VGND VGND VPWR VPWR _21722_/X sky130_fd_sc_hd__o22a_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21653_ _21192_/X _21653_/B _21653_/C VGND VGND VPWR VPWR _21653_/X sky130_fd_sc_hd__and3_4
X_24441_ _24459_/CLK _24441_/D HRESETn VGND VGND VPWR VPWR _22365_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20793__B _20792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20604_ _20598_/X _20600_/Y _24168_/Q _20603_/X VGND VGND VPWR VPWR _23737_/D sky130_fd_sc_hd__a2bb2o_4
X_21584_ _21583_/X VGND VGND VPWR VPWR _22006_/B sky130_fd_sc_hd__buf_2
X_24372_ _24372_/CLK _15971_/X HRESETn VGND VGND VPWR VPWR _15970_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_71_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23831__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20535_ _20534_/Y _20531_/Y _13514_/X VGND VGND VPWR VPWR _20535_/X sky130_fd_sc_hd__o21a_4
X_23323_ _24750_/CLK _19476_/X VGND VGND VPWR VPWR _23323_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25055__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13356__B2 _13338_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20466_ _20465_/X VGND VGND VPWR VPWR _20466_/X sky130_fd_sc_hd__buf_2
X_23254_ _23278_/CLK _19669_/X VGND VGND VPWR VPWR _19665_/A sky130_fd_sc_hd__dfxtp_4
X_22205_ _21175_/X _22202_/X _22203_/X _22205_/D VGND VGND VPWR VPWR _22205_/X sky130_fd_sc_hd__or4_4
X_23185_ _25050_/CLK _19855_/X VGND VGND VPWR VPWR _19853_/A sky130_fd_sc_hd__dfxtp_4
X_20397_ _17183_/A _20394_/A _17184_/Y VGND VGND VPWR VPWR _20397_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22136_ _21245_/X _22133_/X _22136_/C _22136_/D VGND VGND VPWR VPWR _22136_/X sky130_fd_sc_hd__or4_4
XFILLER_121_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14305__B1 _14304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14856__B2 _14835_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22067_ _21396_/A _22059_/X _22066_/X VGND VGND VPWR VPWR _22067_/X sky130_fd_sc_hd__and3_4
XFILLER_59_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19741__A2_N _19738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24690__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21018_ _14469_/X _20997_/Y _21004_/Y _21011_/Y _21017_/Y VGND VGND VPWR VPWR _21018_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_48_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13840_ _13830_/X _13839_/X VGND VGND VPWR VPWR _13840_/Y sky130_fd_sc_hd__nor2_4
XFILLER_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12070__A1_N _20889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19547__B2 _19546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21145__A _21335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13771_ _13771_/A VGND VGND VPWR VPWR _14073_/B sky130_fd_sc_hd__inv_2
XFILLER_74_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19756__A2_N _19750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22969_ _24390_/Q _22834_/B VGND VGND VPWR VPWR _22969_/X sky130_fd_sc_hd__or2_4
X_15510_ _12085_/Y _15509_/X _13658_/X _15509_/X VGND VGND VPWR VPWR _24555_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_69_0_HCLK clkbuf_6_34_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_69_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12722_ _12609_/A _12722_/B VGND VGND VPWR VPWR _12722_/X sky130_fd_sc_hd__or2_4
X_24708_ _24674_/CLK _24708_/D HRESETn VGND VGND VPWR VPWR _24708_/Q sky130_fd_sc_hd__dfrtp_4
X_16490_ _24184_/Q VGND VGND VPWR VPWR _16490_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20984__A _20979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15441_ _15439_/X _15441_/B VGND VGND VPWR VPWR _15452_/B sky130_fd_sc_hd__or2_4
XANTENNA__23919__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12653_ _12731_/A _12728_/A _12653_/C VGND VGND VPWR VPWR _12653_/X sky130_fd_sc_hd__or3_4
XFILLER_31_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24639_ _23762_/CLK _15263_/X HRESETn VGND VGND VPWR VPWR _13728_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21799__B _21181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16781__A1 _15862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ HWDATA[9] VGND VGND VPWR VPWR _11604_/X sky130_fd_sc_hd__buf_2
X_18160_ _16121_/A _18159_/A _16121_/Y _18327_/A VGND VGND VPWR VPWR _18160_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15372_ _22408_/A _15366_/X _11590_/X _15366_/X VGND VGND VPWR VPWR _15372_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _12584_/A VGND VGND VPWR VPWR _12584_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17111_ _17108_/B VGND VGND VPWR VPWR _17112_/B sky130_fd_sc_hd__inv_2
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14323_ _20177_/A _14321_/X _14329_/A _14322_/Y VGND VGND VPWR VPWR _14323_/X sky130_fd_sc_hd__a211o_4
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11535_ _15920_/A VGND VGND VPWR VPWR _11535_/X sky130_fd_sc_hd__buf_2
X_18091_ _21644_/A VGND VGND VPWR VPWR _18091_/Y sky130_fd_sc_hd__inv_2
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17042_ _17042_/A _16992_/Y _16982_/Y _17042_/D VGND VGND VPWR VPWR _17042_/X sky130_fd_sc_hd__or4_4
XANTENNA__12933__C _12933_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14254_ _14252_/Y _14249_/X _14236_/X _14253_/X VGND VGND VPWR VPWR _14254_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13205_ _13301_/A _13205_/B VGND VGND VPWR VPWR _13206_/C sky130_fd_sc_hd__or2_4
X_14185_ _14175_/X _14184_/X _25152_/Q _14180_/X VGND VGND VPWR VPWR _14185_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19483__B1 _19366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16702__A _22782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24778__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13136_ _13136_/A _19333_/A VGND VGND VPWR VPWR _13138_/B sky130_fd_sc_hd__or2_4
XANTENNA__12570__A2 _24510_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18993_ _23493_/Q VGND VGND VPWR VPWR _21940_/B sky130_fd_sc_hd__inv_2
XANTENNA__24707__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14847__B2 _24137_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15318__A _16231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13067_ _13076_/A VGND VGND VPWR VPWR _13300_/A sky130_fd_sc_hd__buf_2
X_17944_ _17944_/A _19075_/A VGND VGND VPWR VPWR _17944_/X sky130_fd_sc_hd__or2_4
XFILLER_117_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16049__B1 _11522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12018_ _12016_/A _12016_/B _12017_/Y VGND VGND VPWR VPWR _12019_/B sky130_fd_sc_hd__o21a_4
X_17875_ _15730_/X _17859_/X _17874_/X _23930_/Q _17765_/X VGND VGND VPWR VPWR _17875_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__21593__A1 _16464_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24360__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22790__B1 _22536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19614_ _19614_/A VGND VGND VPWR VPWR _19614_/X sky130_fd_sc_hd__buf_2
X_16826_ _16765_/Y _16823_/Y _16826_/C _16825_/Y VGND VGND VPWR VPWR _16827_/C sky130_fd_sc_hd__or4_4
XANTENNA__12038__A1_N _11992_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14876__B _15034_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16757_ _15866_/Y _24075_/Q _15866_/Y _24075_/Q VGND VGND VPWR VPWR _16757_/X sky130_fd_sc_hd__a2bb2o_4
X_19545_ _19545_/A VGND VGND VPWR VPWR _21328_/B sky130_fd_sc_hd__inv_2
X_13969_ _24890_/Q _13928_/X _24890_/Q _13928_/X VGND VGND VPWR VPWR _13969_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12677__A _12638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11581__A _16087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15708_ _12349_/Y _15702_/X _15286_/X _15702_/X VGND VGND VPWR VPWR _24469_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15053__A _15019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16688_ _16683_/X _16688_/B _16686_/X _16687_/X VGND VGND VPWR VPWR _16717_/A sky130_fd_sc_hd__or4_4
X_19476_ _19475_/Y _19473_/X _19381_/X _19473_/X VGND VGND VPWR VPWR _19476_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15639_ _21088_/A VGND VGND VPWR VPWR _15639_/X sky130_fd_sc_hd__buf_2
X_18427_ _18427_/A _18427_/B _18427_/C _18426_/X VGND VGND VPWR VPWR _18485_/D sky130_fd_sc_hd__or4_4
XANTENNA__16772__A1 _15889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18358_ _23831_/Q VGND VGND VPWR VPWR _18358_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22845__A1 _23026_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22845__B2 _22460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18083__B _18080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17309_ _17309_/A VGND VGND VPWR VPWR _17382_/C sky130_fd_sc_hd__inv_2
X_18289_ _18289_/A VGND VGND VPWR VPWR _18289_/Y sky130_fd_sc_hd__inv_2
X_20320_ _14255_/Y _20296_/A _20286_/X _20319_/X VGND VGND VPWR VPWR _20320_/X sky130_fd_sc_hd__a211o_4
XFILLER_128_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20251_ _20251_/A _20251_/B VGND VGND VPWR VPWR _20252_/D sky130_fd_sc_hd__and2_4
XANTENNA__19474__B1 _19424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16288__B1 _24259_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20182_ _20189_/A _20181_/X VGND VGND VPWR VPWR _20182_/X sky130_fd_sc_hd__or2_4
XFILLER_118_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24448__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24990_ _24841_/CLK _24990_/D HRESETn VGND VGND VPWR VPWR _13348_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_69_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23941_ _23343_/CLK _23941_/D HRESETn VGND VGND VPWR VPWR _23941_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23872_ _23872_/CLK _23872_/D HRESETn VGND VGND VPWR VPWR _18244_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24030__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18258__B _18459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22823_ _24314_/Q _22897_/B VGND VGND VPWR VPWR _22823_/X sky130_fd_sc_hd__or2_4
XANTENNA__12077__B2 _12089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22754_ _21561_/X _22752_/X _21562_/X _22753_/X VGND VGND VPWR VPWR _22754_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16212__B1 _16211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21705_ _21793_/A _21705_/B _21705_/C VGND VGND VPWR VPWR _21705_/X sky130_fd_sc_hd__and3_4
XFILLER_25_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22685_ _22685_/A VGND VGND VPWR VPWR _22686_/C sky130_fd_sc_hd__inv_2
XFILLER_90_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24424_ _24399_/CLK _15835_/X HRESETn VGND VGND VPWR VPWR _24424_/Q sky130_fd_sc_hd__dfrtp_4
X_21636_ _20745_/X _21620_/X _21635_/X VGND VGND VPWR VPWR _21636_/X sky130_fd_sc_hd__and3_4
XANTENNA__22836__A1 _22335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21639__A2 _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22836__B2 _22576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24355_ _24349_/CLK _24355_/D HRESETn VGND VGND VPWR VPWR _24355_/Q sky130_fd_sc_hd__dfrtp_4
X_21567_ _21567_/A _22445_/B VGND VGND VPWR VPWR _21567_/X sky130_fd_sc_hd__and2_4
XFILLER_21_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23306_ _23282_/CLK _23306_/D VGND VGND VPWR VPWR _19520_/A sky130_fd_sc_hd__dfxtp_4
X_20518_ _23717_/Q _20513_/X _20517_/Y VGND VGND VPWR VPWR _20518_/Y sky130_fd_sc_hd__a21oi_4
X_21498_ _21367_/A _19498_/Y VGND VGND VPWR VPWR _21498_/X sky130_fd_sc_hd__or2_4
XFILLER_14_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24286_ _24138_/CLK _24286_/D HRESETn VGND VGND VPWR VPWR _24286_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20449_ _20448_/X VGND VGND VPWR VPWR _20453_/B sky130_fd_sc_hd__buf_2
XANTENNA__17618__A _17615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19465__B1 _18662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23237_ _23246_/CLK _23237_/D VGND VGND VPWR VPWR _19713_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_10_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21272__B1 _21062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18440__C _18459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23168_ _25112_/CLK _19900_/X VGND VGND VPWR VPWR _19899_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24189__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22119_ _22116_/X _22117_/X _21974_/X _25197_/Q _22118_/X VGND VGND VPWR VPWR _22120_/B
+ sky130_fd_sc_hd__a32o_4
X_15990_ _15989_/Y _15987_/X _15897_/X _15987_/X VGND VGND VPWR VPWR _24365_/D sky130_fd_sc_hd__a2bb2o_4
X_23099_ _23258_/CLK _20083_/X VGND VGND VPWR VPWR _23099_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24118__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20979__A _20979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14941_ _24664_/Q VGND VGND VPWR VPWR _14941_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22367__A3 _21981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17660_ _13406_/A VGND VGND VPWR VPWR _17662_/A sky130_fd_sc_hd__inv_2
X_14872_ _14742_/Y _14872_/B _15078_/A _14871_/X VGND VGND VPWR VPWR _14873_/D sky130_fd_sc_hd__or4_4
XFILLER_76_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16611_ _14836_/Y _16606_/X _16373_/X _16610_/X VGND VGND VPWR VPWR _16611_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22119__A3 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13823_ _24905_/Q VGND VGND VPWR VPWR _13869_/B sky130_fd_sc_hd__inv_2
X_17591_ _22307_/A _17591_/B VGND VGND VPWR VPWR _17591_/X sky130_fd_sc_hd__or2_4
XFILLER_91_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16542_ _16530_/A VGND VGND VPWR VPWR _16542_/X sky130_fd_sc_hd__buf_2
X_19330_ _19325_/Y _19328_/X _19329_/X _19328_/X VGND VGND VPWR VPWR _19330_/X sky130_fd_sc_hd__a2bb2o_4
X_13754_ _13754_/A _13754_/B _13722_/A _24635_/Q VGND VGND VPWR VPWR _13773_/D sky130_fd_sc_hd__or4_4
XFILLER_44_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12705_ _12716_/A _12703_/X _12705_/C VGND VGND VPWR VPWR _25058_/D sky130_fd_sc_hd__and3_4
X_19261_ _19260_/X VGND VGND VPWR VPWR _19261_/X sky130_fd_sc_hd__buf_2
XANTENNA__21603__A _17651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23753__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16473_ _24190_/Q VGND VGND VPWR VPWR _16473_/Y sky130_fd_sc_hd__inv_2
X_13685_ _20201_/A _13683_/X _13678_/X _13684_/Y VGND VGND VPWR VPWR _24923_/D sky130_fd_sc_hd__a211o_4
X_18212_ _18212_/A VGND VGND VPWR VPWR _18212_/Y sky130_fd_sc_hd__inv_2
X_15424_ _12062_/A VGND VGND VPWR VPWR _15424_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12636_ _12963_/A VGND VGND VPWR VPWR _12636_/X sky130_fd_sc_hd__buf_2
X_19192_ _19188_/Y _19191_/X _19170_/X _19191_/X VGND VGND VPWR VPWR _19192_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_156_0_HCLK clkbuf_7_78_0_HCLK/X VGND VGND VPWR VPWR _24435_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18143_ _24345_/Q _18268_/A _16056_/A _18221_/A VGND VGND VPWR VPWR _18145_/C sky130_fd_sc_hd__a2bb2o_4
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15355_ _24603_/Q VGND VGND VPWR VPWR _22624_/A sky130_fd_sc_hd__inv_2
X_12567_ _25056_/Q _24521_/Q _12565_/Y _12566_/Y VGND VGND VPWR VPWR _12577_/A sky130_fd_sc_hd__o22a_4
XFILLER_129_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24959__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14306_ _14306_/A VGND VGND VPWR VPWR _14306_/Y sky130_fd_sc_hd__inv_2
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11518_ _11537_/A VGND VGND VPWR VPWR _11518_/Y sky130_fd_sc_hd__inv_2
X_18074_ _11755_/A VGND VGND VPWR VPWR _19303_/A sky130_fd_sc_hd__buf_2
X_15286_ _15801_/A VGND VGND VPWR VPWR _15286_/X sky130_fd_sc_hd__buf_2
X_12498_ _12498_/A _12495_/X VGND VGND VPWR VPWR _12499_/C sky130_fd_sc_hd__or2_4
XANTENNA__22434__A _22434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23664__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17025_ _17080_/A VGND VGND VPWR VPWR _17026_/A sky130_fd_sc_hd__inv_2
X_14237_ _14226_/A VGND VGND VPWR VPWR _14237_/X sky130_fd_sc_hd__buf_2
XANTENNA__22153__B _22153_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14168_ _14168_/A VGND VGND VPWR VPWR _14169_/B sky130_fd_sc_hd__inv_2
XANTENNA__24541__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11576__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13119_ _13297_/A _23556_/Q VGND VGND VPWR VPWR _13119_/X sky130_fd_sc_hd__or2_4
XANTENNA__19208__B1 _19207_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14099_ _14099_/A VGND VGND VPWR VPWR _15260_/A sky130_fd_sc_hd__buf_2
X_18976_ _18974_/Y _18970_/X _18883_/X _18975_/X VGND VGND VPWR VPWR _18976_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20889__A _20889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17927_ _17927_/A _19094_/A VGND VGND VPWR VPWR _17929_/B sky130_fd_sc_hd__or2_4
XFILLER_38_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17858_ _17738_/A _17858_/B _17857_/X VGND VGND VPWR VPWR _17859_/C sky130_fd_sc_hd__or3_4
XFILLER_82_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16442__B1 _16093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16809_ _16809_/A _16806_/X _16809_/C _16808_/X VGND VGND VPWR VPWR _16810_/D sky130_fd_sc_hd__or4_4
XFILLER_93_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17789_ _17894_/A _17789_/B _17788_/X VGND VGND VPWR VPWR _17794_/B sky130_fd_sc_hd__and3_4
XFILLER_81_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19528_ _19527_/Y _19523_/X _19506_/X _19510_/Y VGND VGND VPWR VPWR _19528_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21869__A2 _20819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_52_0_HCLK clkbuf_6_26_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_52_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19459_ _15556_/X VGND VGND VPWR VPWR _19459_/X sky130_fd_sc_hd__buf_2
XANTENNA__15511__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22470_ _13360_/A _22469_/X _21058_/X _24560_/Q _21059_/X VGND VGND VPWR VPWR _22470_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22818__B2 _21187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21421_ _16381_/A _21553_/A _21292_/X _21420_/X VGND VGND VPWR VPWR _21422_/C sky130_fd_sc_hd__a211o_4
XFILLER_136_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21352_ _21352_/A _21352_/B VGND VGND VPWR VPWR _21353_/C sky130_fd_sc_hd__or2_4
X_24140_ _24140_/CLK _16596_/X HRESETn VGND VGND VPWR VPWR _16594_/A sky130_fd_sc_hd__dfrtp_4
X_20303_ _18614_/B _20301_/Y _20315_/C VGND VGND VPWR VPWR _20303_/X sky130_fd_sc_hd__and3_4
XFILLER_50_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21283_ _21867_/A VGND VGND VPWR VPWR _22407_/A sky130_fd_sc_hd__buf_2
X_24071_ _24071_/CLK _24071_/D HRESETn VGND VGND VPWR VPWR _24071_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20234_ _13891_/A _20234_/B VGND VGND VPWR VPWR _20234_/X sky130_fd_sc_hd__and2_4
X_23022_ _16304_/A _15919_/X _22858_/X _23021_/X VGND VGND VPWR VPWR _23022_/X sky130_fd_sc_hd__a211o_4
XFILLER_89_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24282__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20165_ _20165_/A VGND VGND VPWR VPWR _20165_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20799__A _22148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24211__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16681__B1 _13463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20096_ _20034_/A _19644_/X _19236_/X VGND VGND VPWR VPWR _20097_/A sky130_fd_sc_hd__or3_4
X_24973_ _24974_/CLK _24973_/D HRESETn VGND VGND VPWR VPWR _24973_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22754__B1 _21562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21557__B2 _21400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22510__C _22510_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23924_ _25159_/CLK _23924_/D HRESETn VGND VGND VPWR VPWR _22450_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21407__B _21324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23855_ _24879_/CLK _23855_/D HRESETn VGND VGND VPWR VPWR _23855_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22506__B1 _22351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17901__A _17716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22806_ _24215_/Q _22806_/B VGND VGND VPWR VPWR _22806_/X sky130_fd_sc_hd__or2_4
X_23786_ _23789_/CLK _23786_/D HRESETn VGND VGND VPWR VPWR _11883_/A sky130_fd_sc_hd__dfrtp_4
X_20998_ _20998_/A _20998_/B VGND VGND VPWR VPWR _21000_/B sky130_fd_sc_hd__or2_4
XFILLER_77_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22737_ _24567_/Q _22557_/X _22558_/X _22736_/X VGND VGND VPWR VPWR _22738_/C sky130_fd_sc_hd__a211o_4
XANTENNA__25070__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16736__B2 _17497_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16517__A _24173_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15421__A _16228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13470_ _13464_/X _13470_/B VGND VGND VPWR VPWR _13475_/A sky130_fd_sc_hd__and2_4
XFILLER_125_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22668_ _21529_/X _22666_/X _13362_/A _22667_/X VGND VGND VPWR VPWR _22668_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_8_229_0_HCLK clkbuf_8_229_0_HCLK/A VGND VGND VPWR VPWR _24185_/CLK sky130_fd_sc_hd__clkbuf_1
X_12421_ _12305_/Y _12419_/A VGND VGND VPWR VPWR _12421_/X sky130_fd_sc_hd__or2_4
X_24407_ _24412_/CLK _24407_/D HRESETn VGND VGND VPWR VPWR _24407_/Q sky130_fd_sc_hd__dfrtp_4
X_21619_ _21614_/X _21618_/X _17639_/A VGND VGND VPWR VPWR _21619_/X sky130_fd_sc_hd__o21a_4
XFILLER_16_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22599_ _22369_/X _22598_/X _21986_/X _11568_/A _21987_/X VGND VGND VPWR VPWR _22599_/X
+ sky130_fd_sc_hd__a32o_4
X_15140_ _24677_/Q _15144_/B VGND VGND VPWR VPWR _15140_/X sky130_fd_sc_hd__or2_4
X_12352_ _12312_/X _12352_/B _12337_/X _12352_/D VGND VGND VPWR VPWR _12398_/A sky130_fd_sc_hd__or4_4
X_24338_ _24349_/CLK _24338_/D HRESETn VGND VGND VPWR VPWR _24338_/Q sky130_fd_sc_hd__dfrtp_4
X_15071_ _15067_/B _15071_/B VGND VGND VPWR VPWR _15075_/B sky130_fd_sc_hd__or2_4
XANTENNA__17348__A _17303_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12283_ _12157_/Y _12283_/B VGND VGND VPWR VPWR _12285_/B sky130_fd_sc_hd__nand2_4
X_24269_ _24140_/CLK _24269_/D HRESETn VGND VGND VPWR VPWR _24269_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15711__A2 _15460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14022_ _14197_/A _14046_/A VGND VGND VPWR VPWR _14037_/B sky130_fd_sc_hd__or2_4
XFILLER_49_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18830_ _23550_/Q VGND VGND VPWR VPWR _22053_/B sky130_fd_sc_hd__inv_2
XFILLER_84_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16672__B1 _16671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15973_ _15987_/A VGND VGND VPWR VPWR _15973_/X sky130_fd_sc_hd__buf_2
X_18761_ _18734_/D _19100_/A VGND VGND VPWR VPWR _18776_/A sky130_fd_sc_hd__nor2_4
XANTENNA__20502__A _13509_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14924_ _24659_/Q _24264_/Q _15208_/A _14923_/Y VGND VGND VPWR VPWR _14924_/X sky130_fd_sc_hd__o22a_4
X_17712_ _17916_/A _17712_/B VGND VGND VPWR VPWR _17715_/B sky130_fd_sc_hd__or2_4
X_18692_ _18697_/A VGND VGND VPWR VPWR _18692_/X sky130_fd_sc_hd__buf_2
XFILLER_75_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16424__B1 _16259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23934__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14855_ _14849_/X _14855_/B _14855_/C _14855_/D VGND VGND VPWR VPWR _14855_/X sky130_fd_sc_hd__or4_4
X_17643_ _17642_/Y VGND VGND VPWR VPWR _17644_/A sky130_fd_sc_hd__buf_2
XANTENNA__25158__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20771__A2 _22201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13806_ _24902_/Q VGND VGND VPWR VPWR _13806_/X sky130_fd_sc_hd__buf_2
XANTENNA__13116__A _13054_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17811__A _17727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17574_ _17547_/X _17572_/X _17573_/X VGND VGND VPWR VPWR _23957_/D sky130_fd_sc_hd__and3_4
X_14786_ _14870_/A _24096_/Q _24683_/Q _14754_/Y VGND VGND VPWR VPWR _14786_/X sky130_fd_sc_hd__a2bb2o_4
X_11998_ _11997_/Y _11995_/X _11616_/X _11995_/X VGND VGND VPWR VPWR _11998_/X sky130_fd_sc_hd__a2bb2o_4
X_16525_ _24170_/Q VGND VGND VPWR VPWR _22343_/A sky130_fd_sc_hd__inv_2
X_19313_ _19310_/Y _19305_/X _19311_/X _19312_/X VGND VGND VPWR VPWR _23380_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21333__A _21333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13737_ _13737_/A VGND VGND VPWR VPWR _13737_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_39_0_HCLK clkbuf_6_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_78_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16727__B2 _22395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16456_ _16454_/Y _16452_/X _16455_/X _16452_/X VGND VGND VPWR VPWR _16456_/X sky130_fd_sc_hd__a2bb2o_4
X_19244_ _19238_/Y VGND VGND VPWR VPWR _19244_/X sky130_fd_sc_hd__buf_2
X_13668_ _13668_/A VGND VGND VPWR VPWR _13668_/X sky130_fd_sc_hd__buf_2
X_15407_ _15407_/A VGND VGND VPWR VPWR _15407_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12619_ _12619_/A VGND VGND VPWR VPWR _12619_/Y sky130_fd_sc_hd__inv_2
X_19175_ _19175_/A VGND VGND VPWR VPWR _19175_/X sky130_fd_sc_hd__buf_2
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16387_ _24222_/Q VGND VGND VPWR VPWR _16387_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13599_ _13558_/B _13598_/Y _13594_/X _13586_/X _11650_/A VGND VGND VPWR VPWR _24951_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24793__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18126_ _18124_/Y _18125_/X _18127_/A _18125_/X VGND VGND VPWR VPWR _18126_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15338_ _15337_/Y _15333_/X _11545_/X _15333_/X VGND VGND VPWR VPWR _15338_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24722__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11972__B1 _11620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18057_ _18045_/X VGND VGND VPWR VPWR _18060_/A sky130_fd_sc_hd__inv_2
XFILLER_117_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15269_ _14100_/X _23767_/Q _15251_/Y _13742_/C _15251_/B VGND VGND VPWR VPWR _24633_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17008_ _24047_/Q VGND VGND VPWR VPWR _17097_/A sky130_fd_sc_hd__inv_2
XFILLER_126_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20039__B2 _20036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21508__A _21214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18959_ _16291_/A VGND VGND VPWR VPWR _18959_/X sky130_fd_sc_hd__buf_2
X_21970_ _21256_/X VGND VGND VPWR VPWR _22306_/A sky130_fd_sc_hd__buf_2
XFILLER_66_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16415__B1 _16251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23675__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20921_ _22445_/B VGND VGND VPWR VPWR _21553_/A sky130_fd_sc_hd__buf_2
XFILLER_81_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20762__A2 _14015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13026__A _13271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17721__A _17721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23640_ _24811_/CLK _23640_/D HRESETn VGND VGND VPWR VPWR _23640_/Q sky130_fd_sc_hd__dfrtp_4
X_20852_ _20852_/A _20852_/B VGND VGND VPWR VPWR _20852_/Y sky130_fd_sc_hd__nor2_4
XPHY_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23571_ _23560_/CLK _23571_/D VGND VGND VPWR VPWR _18771_/A sky130_fd_sc_hd__dfxtp_4
X_20783_ _20751_/X VGND VGND VPWR VPWR _20783_/X sky130_fd_sc_hd__buf_2
XANTENNA__21711__A1 _15322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21711__B2 _22148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22522_ _22369_/X _22521_/X _21986_/X _11575_/A _21987_/X VGND VGND VPWR VPWR _22522_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16785__A1_N _24412_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22453_ _20617_/Y _21576_/X _20480_/Y _22452_/X VGND VGND VPWR VPWR _22453_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13401__B1 _13330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21404_ _22146_/B _21401_/X _21256_/X _21403_/X VGND VGND VPWR VPWR _21404_/X sky130_fd_sc_hd__a211o_4
XFILLER_136_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25172_ _23246_/CLK _11849_/X HRESETn VGND VGND VPWR VPWR _19724_/A sky130_fd_sc_hd__dfrtp_4
X_22384_ _21991_/X _22383_/X VGND VGND VPWR VPWR _22384_/X sky130_fd_sc_hd__and2_4
XANTENNA__24463__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_59_0_HCLK clkbuf_8_59_0_HCLK/A VGND VGND VPWR VPWR _25217_/CLK sky130_fd_sc_hd__clkbuf_1
X_24123_ _24698_/CLK _16626_/X HRESETn VGND VGND VPWR VPWR _24123_/Q sky130_fd_sc_hd__dfrtp_4
X_21335_ _21335_/A _21335_/B VGND VGND VPWR VPWR _21337_/B sky130_fd_sc_hd__or2_4
XFILLER_136_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24054_ _24612_/CLK _17071_/X HRESETn VGND VGND VPWR VPWR _24054_/Q sky130_fd_sc_hd__dfrtp_4
X_21266_ _24362_/Q _21043_/X VGND VGND VPWR VPWR _21266_/X sky130_fd_sc_hd__or2_4
XANTENNA__22802__A _24118_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23005_ _24460_/Q _22015_/X VGND VGND VPWR VPWR _23005_/X sky130_fd_sc_hd__or2_4
X_20217_ _23690_/Q VGND VGND VPWR VPWR _20217_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16249__A3 _15477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21197_ _21367_/A _21197_/B VGND VGND VPWR VPWR _21201_/B sky130_fd_sc_hd__or2_4
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16654__B1 _24107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20148_ _20141_/A VGND VGND VPWR VPWR _20148_/X sky130_fd_sc_hd__buf_2
XANTENNA__20322__A _24805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22727__B1 _14960_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11944__A _22477_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15416__A _13644_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12970_ _12969_/X VGND VGND VPWR VPWR _25017_/D sky130_fd_sc_hd__inv_2
X_20079_ _23100_/Q VGND VGND VPWR VPWR _21909_/B sky130_fd_sc_hd__inv_2
XANTENNA__19650__A1_N _21935_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24956_ _24757_/CLK _13588_/X HRESETn VGND VGND VPWR VPWR _11685_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_44_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11921_ _25163_/Q VGND VGND VPWR VPWR _21897_/A sky130_fd_sc_hd__inv_2
X_23907_ _23908_/CLK _23907_/D HRESETn VGND VGND VPWR VPWR _18011_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_73_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24887_ _23774_/CLK _13982_/X HRESETn VGND VGND VPWR VPWR _24887_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14640_ _14620_/Y VGND VGND VPWR VPWR _14640_/X sky130_fd_sc_hd__buf_2
XFILLER_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11852_ _11830_/Y VGND VGND VPWR VPWR _11852_/X sky130_fd_sc_hd__buf_2
X_23838_ _23828_/CLK _23838_/D HRESETn VGND VGND VPWR VPWR _23838_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15364__A1_N _15363_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22249__A _22249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21153__A _21153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14571_ _17742_/A VGND VGND VPWR VPWR _14571_/X sky130_fd_sc_hd__buf_2
X_11783_ _11809_/A _11782_/X VGND VGND VPWR VPWR _11783_/X sky130_fd_sc_hd__or2_4
XANTENNA__13640__B1 _13638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23769_ _24728_/CLK _23769_/D HRESETn VGND VGND VPWR VPWR _20244_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20505__A2 _20416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16310_ _16310_/A VGND VGND VPWR VPWR _16310_/Y sky130_fd_sc_hd__inv_2
X_13522_ _24965_/Q _13388_/X _13521_/Y VGND VGND VPWR VPWR _24965_/D sky130_fd_sc_hd__o21a_4
XFILLER_57_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17290_ _17283_/X _17290_/B _17290_/C _17289_/X VGND VGND VPWR VPWR _17296_/C sky130_fd_sc_hd__or4_4
XFILLER_9_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16241_ _16256_/A VGND VGND VPWR VPWR _16247_/A sky130_fd_sc_hd__buf_2
X_13453_ _13443_/X _13453_/B _13448_/X _13453_/D VGND VGND VPWR VPWR _13453_/X sky130_fd_sc_hd__or4_4
XFILLER_51_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14990__A _14990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12404_ _21104_/A VGND VGND VPWR VPWR _12536_/A sky130_fd_sc_hd__inv_2
X_16172_ _16172_/A VGND VGND VPWR VPWR _16172_/Y sky130_fd_sc_hd__inv_2
X_13384_ _20691_/B VGND VGND VPWR VPWR _20688_/B sky130_fd_sc_hd__buf_2
XANTENNA__21600__B _21600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15123_ _15123_/A _15123_/B VGND VGND VPWR VPWR _15123_/X sky130_fd_sc_hd__and2_4
XFILLER_5_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12335_ _24474_/Q VGND VGND VPWR VPWR _12335_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24133__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15054_ _15018_/X _15052_/X _15054_/C VGND VGND VPWR VPWR _15054_/X sky130_fd_sc_hd__and3_4
X_19931_ _23156_/Q VGND VGND VPWR VPWR _21766_/B sky130_fd_sc_hd__inv_2
XFILLER_126_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12266_ _12180_/B _12265_/X VGND VGND VPWR VPWR _12267_/B sky130_fd_sc_hd__or2_4
XFILLER_107_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22712__A _22712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14005_ _13925_/B _14000_/B _14000_/Y VGND VGND VPWR VPWR _14005_/Y sky130_fd_sc_hd__a21oi_4
X_19862_ _19862_/A _19862_/B _19883_/C VGND VGND VPWR VPWR _19863_/A sky130_fd_sc_hd__or3_4
X_12197_ _12196_/X VGND VGND VPWR VPWR _12197_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16645__B1 _16264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22431__B _22505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18813_ _23556_/Q VGND VGND VPWR VPWR _18813_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19793_ _19780_/Y VGND VGND VPWR VPWR _19793_/X sky130_fd_sc_hd__buf_2
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15326__A _15401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18744_ _18743_/X VGND VGND VPWR VPWR _18744_/X sky130_fd_sc_hd__buf_2
X_15956_ _15955_/Y _15953_/X _15775_/X _15953_/X VGND VGND VPWR VPWR _15956_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14907_ _24274_/Q VGND VGND VPWR VPWR _14907_/Y sky130_fd_sc_hd__inv_2
X_15887_ _24403_/Q VGND VGND VPWR VPWR _15887_/Y sky130_fd_sc_hd__inv_2
X_18675_ _23603_/Q VGND VGND VPWR VPWR _18675_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20886__B _11725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17626_ _17459_/Y _17625_/Y _17447_/Y VGND VGND VPWR VPWR _17626_/X sky130_fd_sc_hd__o21a_4
X_14838_ _24142_/Q VGND VGND VPWR VPWR _14838_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15620__A1 _15619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22159__A _11961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15620__B2 _15585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14769_ _15034_/A _14751_/A _14712_/X _14713_/Y VGND VGND VPWR VPWR _14769_/X sky130_fd_sc_hd__a2bb2o_4
X_17557_ _17556_/X VGND VGND VPWR VPWR _23962_/D sky130_fd_sc_hd__inv_2
XANTENNA__19898__B1 _19832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24974__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16508_ _24177_/Q VGND VGND VPWR VPWR _16508_/Y sky130_fd_sc_hd__inv_2
X_17488_ _20778_/A VGND VGND VPWR VPWR _17488_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24903__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19227_ _11635_/A VGND VGND VPWR VPWR _19227_/X sky130_fd_sc_hd__buf_2
XFILLER_108_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16439_ _16452_/A VGND VGND VPWR VPWR _16439_/X sky130_fd_sc_hd__buf_2
XFILLER_34_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15384__B1 _11607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_212_0_HCLK clkbuf_8_213_0_HCLK/A VGND VGND VPWR VPWR _24192_/CLK sky130_fd_sc_hd__clkbuf_1
X_19158_ _19157_/Y _19153_/X _19089_/X _19153_/X VGND VGND VPWR VPWR _19158_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18109_ _18108_/Y _18096_/Y _18093_/A _18095_/X VGND VGND VPWR VPWR _23886_/D sky130_fd_sc_hd__o22a_4
XFILLER_121_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19089_ _18678_/X VGND VGND VPWR VPWR _19089_/X sky130_fd_sc_hd__buf_2
X_21120_ SSn_S2 _13324_/X VGND VGND VPWR VPWR _21120_/X sky130_fd_sc_hd__or2_4
XFILLER_132_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21051_ _21050_/Y VGND VGND VPWR VPWR _21051_/X sky130_fd_sc_hd__buf_2
XFILLER_132_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22421__A2 _20799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20002_ _23129_/Q VGND VGND VPWR VPWR _20002_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12370__B1 _12415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16636__B1 HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23856__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24810_ _24788_/CLK _24810_/D HRESETn VGND VGND VPWR VPWR _24810_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__22185__A1 _22155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25009__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22185__B2 _22884_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24741_ _24740_/CLK _14547_/X HRESETn VGND VGND VPWR VPWR _24741_/Q sky130_fd_sc_hd__dfrtp_4
X_21953_ _21214_/A _21953_/B VGND VGND VPWR VPWR _21955_/B sky130_fd_sc_hd__or2_4
XFILLER_27_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20904_ _20072_/A _20826_/X _23078_/Q _20827_/X VGND VGND VPWR VPWR _20904_/X sky130_fd_sc_hd__o22a_4
X_24672_ _24676_/CLK _24672_/D HRESETn VGND VGND VPWR VPWR _24672_/Q sky130_fd_sc_hd__dfrtp_4
X_21884_ _21884_/A _22006_/B VGND VGND VPWR VPWR _21884_/Y sky130_fd_sc_hd__nor2_4
XPHY_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ _24769_/CLK _20710_/X HRESETn VGND VGND VPWR VPWR _23623_/Q sky130_fd_sc_hd__dfrtp_4
X_20835_ _16305_/A _20831_/X _20833_/X _20834_/Y VGND VGND VPWR VPWR _20835_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16094__A1_N _22401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_22_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23554_ _23133_/CLK _18820_/X VGND VGND VPWR VPWR _13194_/B sky130_fd_sc_hd__dfxtp_4
X_20766_ _21092_/B VGND VGND VPWR VPWR _20931_/A sky130_fd_sc_hd__buf_2
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24644__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22505_ _22505_/A VGND VGND VPWR VPWR _22505_/X sky130_fd_sc_hd__buf_2
XFILLER_126_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15375__B1 _11594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19378__A _19372_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15914__A2 _15410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23485_ _23482_/CLK _23485_/D VGND VGND VPWR VPWR _23485_/Q sky130_fd_sc_hd__dfxtp_4
X_20697_ _12019_/B _20697_/B VGND VGND VPWR VPWR _20697_/X sky130_fd_sc_hd__and2_4
XFILLER_13_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22436_ _22436_/A _22445_/B VGND VGND VPWR VPWR _22436_/X sky130_fd_sc_hd__and2_4
XFILLER_104_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15127__B1 _15126_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25155_ _24953_/CLK _25155_/D HRESETn VGND VGND VPWR VPWR _25155_/Q sky130_fd_sc_hd__dfrtp_4
X_22367_ _22364_/X _22365_/X _21981_/X _24514_/Q _22366_/X VGND VGND VPWR VPWR _22367_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_109_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12120_ _12120_/A _12093_/X _12106_/X _12119_/X VGND VGND VPWR VPWR _12120_/X sky130_fd_sc_hd__or4_4
X_24106_ _24113_/CLK _24106_/D HRESETn VGND VGND VPWR VPWR _16655_/A sky130_fd_sc_hd__dfrtp_4
X_21318_ _21318_/A VGND VGND VPWR VPWR _21318_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25086_ _25091_/CLK _12485_/Y HRESETn VGND VGND VPWR VPWR _12313_/A sky130_fd_sc_hd__dfrtp_4
X_22298_ _21248_/X _22297_/X _21036_/X _24513_/Q _20780_/A VGND VGND VPWR VPWR _22298_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_117_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12361__A1_N _12495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22948__B1 _14920_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12051_ _12051_/A _20693_/B VGND VGND VPWR VPWR _12051_/X sky130_fd_sc_hd__and2_4
X_24037_ _24037_/CLK _17143_/Y HRESETn VGND VGND VPWR VPWR _16966_/A sky130_fd_sc_hd__dfrtp_4
X_21249_ _21248_/X VGND VGND VPWR VPWR _22146_/B sky130_fd_sc_hd__buf_2
XANTENNA__22412__A2 _22173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16530__A _16530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15810_ _13473_/A _15810_/B VGND VGND VPWR VPWR _15810_/X sky130_fd_sc_hd__and2_4
X_16790_ _15872_/Y _16825_/A _15872_/Y _16825_/A VGND VGND VPWR VPWR _16790_/X sky130_fd_sc_hd__a2bb2o_4
X_15741_ _11944_/X _15741_/B VGND VGND VPWR VPWR _15741_/X sky130_fd_sc_hd__or2_4
XFILLER_86_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12953_ _12943_/C _12943_/D _12922_/X _12951_/B VGND VGND VPWR VPWR _12953_/X sky130_fd_sc_hd__a211o_4
X_24939_ _24937_/CLK _24939_/D HRESETn VGND VGND VPWR VPWR _24939_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_104_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_104_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_11904_ _11904_/A VGND VGND VPWR VPWR _11904_/Y sky130_fd_sc_hd__inv_2
X_15672_ _15689_/A VGND VGND VPWR VPWR _15672_/X sky130_fd_sc_hd__buf_2
X_18460_ _18460_/A VGND VGND VPWR VPWR _18466_/B sky130_fd_sc_hd__inv_2
X_12884_ _12838_/Y _12845_/Y _12884_/C _12883_/X VGND VGND VPWR VPWR _12884_/X sky130_fd_sc_hd__or4_4
X_14623_ _14614_/C VGND VGND VPWR VPWR _14630_/A sky130_fd_sc_hd__inv_2
X_17411_ _17317_/D _17411_/B VGND VGND VPWR VPWR _17412_/B sky130_fd_sc_hd__or2_4
X_11835_ _19597_/A VGND VGND VPWR VPWR _11835_/X sky130_fd_sc_hd__buf_2
X_18391_ _18430_/A VGND VGND VPWR VPWR _18509_/A sky130_fd_sc_hd__buf_2
XFILLER_33_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _24007_/Q _17342_/B VGND VGND VPWR VPWR _17344_/B sky130_fd_sc_hd__or2_4
XPHY_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14553_/Y VGND VGND VPWR VPWR _16035_/B sky130_fd_sc_hd__buf_2
XFILLER_14_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11766_ _11765_/X VGND VGND VPWR VPWR _11766_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14940__A2_N _24267_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24385__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _21887_/A _13505_/B VGND VGND VPWR VPWR _13506_/B sky130_fd_sc_hd__or2_4
X_17273_ _17430_/A VGND VGND VPWR VPWR _17273_/Y sky130_fd_sc_hd__inv_2
XPHY_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ _24745_/Q VGND VGND VPWR VPWR _14485_/Y sky130_fd_sc_hd__inv_2
XPHY_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11697_ _11718_/B VGND VGND VPWR VPWR _11697_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24314__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16224_ _15443_/B _16221_/X _16223_/Y _16224_/D VGND VGND VPWR VPWR _16224_/X sky130_fd_sc_hd__or4_4
X_19012_ _19012_/A VGND VGND VPWR VPWR _19012_/Y sky130_fd_sc_hd__inv_2
X_13436_ _24932_/Q _13435_/A _13434_/Y _13435_/Y VGND VGND VPWR VPWR _13436_/X sky130_fd_sc_hd__o22a_4
XFILLER_70_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_0_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16155_ _24314_/Q VGND VGND VPWR VPWR _16155_/Y sky130_fd_sc_hd__inv_2
X_13367_ _22006_/A _13363_/X _11612_/X _13366_/X VGND VGND VPWR VPWR _13367_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14225__A _14047_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15106_ _15106_/A _15177_/A _15105_/X VGND VGND VPWR VPWR _15107_/C sky130_fd_sc_hd__or3_4
X_12318_ _25080_/Q _12316_/Y _12416_/A _24493_/Q VGND VGND VPWR VPWR _12324_/B sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_42_0_HCLK clkbuf_8_43_0_HCLK/A VGND VGND VPWR VPWR _23531_/CLK sky130_fd_sc_hd__clkbuf_1
X_16086_ _24339_/Q VGND VGND VPWR VPWR _22479_/A sky130_fd_sc_hd__inv_2
X_13298_ _13202_/A _23591_/Q VGND VGND VPWR VPWR _13298_/X sky130_fd_sc_hd__or2_4
X_15037_ _15034_/B VGND VGND VPWR VPWR _15038_/B sky130_fd_sc_hd__inv_2
X_19914_ _21677_/B _19911_/X _19825_/X _19911_/X VGND VGND VPWR VPWR _23163_/D sky130_fd_sc_hd__a2bb2o_4
X_12249_ _12227_/X _12243_/B _12249_/C VGND VGND VPWR VPWR _25118_/D sky130_fd_sc_hd__and3_4
XANTENNA__17536__A _17482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22161__B _22953_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16618__B1 _16617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14879__B _15003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19845_ _21950_/B _19842_/X _19818_/X _19842_/X VGND VGND VPWR VPWR _23189_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25173__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16094__B2 _16090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17291__B1 _25191_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11584__A HWDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19776_ _19776_/A VGND VGND VPWR VPWR _19776_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25102__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16988_ _21291_/A VGND VGND VPWR VPWR _17161_/A sky130_fd_sc_hd__inv_2
XFILLER_37_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18727_ _18726_/Y _18724_/X _18706_/X _18724_/X VGND VGND VPWR VPWR _23585_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15939_ _15938_/Y _15936_/X _11548_/X _15936_/X VGND VGND VPWR VPWR _15939_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18367__A _18359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18658_ _21377_/B _18657_/X _15563_/X _18657_/X VGND VGND VPWR VPWR _23609_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17609_ _23947_/Q _17609_/B VGND VGND VPWR VPWR _17609_/X sky130_fd_sc_hd__or2_4
XFILLER_52_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18589_ _16338_/Y _23832_/Q _16338_/Y _23832_/Q VGND VGND VPWR VPWR _18592_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20620_ _20598_/X _20619_/X _16520_/A _20603_/X VGND VGND VPWR VPWR _20620_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20551_ _20554_/A _20551_/B VGND VGND VPWR VPWR _20601_/A sky130_fd_sc_hd__or2_4
XFILLER_138_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24055__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22336__B _22574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23270_ _23278_/CLK _23270_/D VGND VGND VPWR VPWR _23270_/Q sky130_fd_sc_hd__dfxtp_4
X_20482_ _20480_/Y _20477_/Y _20481_/X VGND VGND VPWR VPWR _20482_/X sky130_fd_sc_hd__o21a_4
XFILLER_20_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22221_ _22216_/X _22354_/A _21246_/X _22220_/X VGND VGND VPWR VPWR _22221_/X sky130_fd_sc_hd__o22a_4
XFILLER_121_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22152_ _22879_/A _22146_/X _22150_/X _15430_/A _22151_/X VGND VGND VPWR VPWR _22183_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_69_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21103_ _21103_/A VGND VGND VPWR VPWR _21128_/C sky130_fd_sc_hd__inv_2
XFILLER_47_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22083_ _11532_/A _20918_/X _22067_/X _22082_/X VGND VGND VPWR VPWR _22083_/X sky130_fd_sc_hd__or4_4
XFILLER_133_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16609__B1 _16369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23690__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21034_ _21033_/X VGND VGND VPWR VPWR _21034_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19810__A3 _13398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22985_ _24155_/Q _22505_/A _22840_/X _22984_/X VGND VGND VPWR VPWR _22986_/C sky130_fd_sc_hd__a211o_4
XANTENNA__24896__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24724_ _24723_/CLK _24724_/D HRESETn VGND VGND VPWR VPWR _14612_/C sky130_fd_sc_hd__dfrtp_4
X_21936_ _21346_/A _21934_/X _21936_/C VGND VGND VPWR VPWR _21936_/X sky130_fd_sc_hd__and3_4
XFILLER_55_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24825__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24655_ _24662_/CLK _24655_/D HRESETn VGND VGND VPWR VPWR _15218_/A sky130_fd_sc_hd__dfrtp_4
X_21867_ _21867_/A VGND VGND VPWR VPWR _22584_/A sky130_fd_sc_hd__buf_2
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _13668_/A VGND VGND VPWR VPWR _11620_/X sky130_fd_sc_hd__buf_2
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ _23990_/CLK _23606_/D VGND VGND VPWR VPWR _23606_/Q sky130_fd_sc_hd__dfxtp_4
X_20818_ _20818_/A VGND VGND VPWR VPWR _20818_/X sky130_fd_sc_hd__buf_2
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24586_ _24013_/CLK _24586_/D HRESETn VGND VGND VPWR VPWR _24586_/Q sky130_fd_sc_hd__dfrtp_4
X_21798_ _23915_/Q _20823_/X _21868_/B _21797_/Y VGND VGND VPWR VPWR _21798_/X sky130_fd_sc_hd__a211o_4
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _11541_/X VGND VGND VPWR VPWR _11551_/X sky130_fd_sc_hd__buf_2
XANTENNA__15348__B1 _11558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23537_ _23537_/CLK _18867_/X VGND VGND VPWR VPWR _13227_/B sky130_fd_sc_hd__dfxtp_4
X_20749_ _20818_/A VGND VGND VPWR VPWR _20749_/X sky130_fd_sc_hd__buf_2
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22246__B _22246_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12128__A2_N _24557_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ _14270_/A VGND VGND VPWR VPWR _14270_/Y sky130_fd_sc_hd__inv_2
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23468_ _23416_/CLK _23468_/D VGND VGND VPWR VPWR _17774_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16560__A2 _16276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13221_ _13221_/A _13219_/X _13221_/C VGND VGND VPWR VPWR _13222_/C sky130_fd_sc_hd__and3_4
XFILLER_137_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25207_ _25012_/CLK _25207_/D HRESETn VGND VGND VPWR VPWR _25207_/Q sky130_fd_sc_hd__dfrtp_4
X_22419_ _22419_/A _11964_/A VGND VGND VPWR VPWR _22419_/X sky130_fd_sc_hd__or2_4
XFILLER_87_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23399_ _23383_/CLK _19257_/X VGND VGND VPWR VPWR _19255_/A sky130_fd_sc_hd__dfxtp_4
X_13152_ _13113_/A _13143_/X _13151_/X VGND VGND VPWR VPWR _13152_/X sky130_fd_sc_hd__and3_4
XFILLER_109_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23778__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_1_0_HCLK clkbuf_8_1_0_HCLK/A VGND VGND VPWR VPWR _23278_/CLK sky130_fd_sc_hd__clkbuf_1
X_25138_ _24980_/CLK _12012_/X HRESETn VGND VGND VPWR VPWR _12011_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_29_0_HCLK clkbuf_6_14_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__22262__A _14047_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12103_ _25109_/Q VGND VGND VPWR VPWR _12103_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23707__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13083_ _13204_/A _18670_/A VGND VGND VPWR VPWR _13083_/X sky130_fd_sc_hd__or2_4
X_17960_ _17928_/A _18756_/A VGND VGND VPWR VPWR _17960_/X sky130_fd_sc_hd__or2_4
X_25069_ _24071_/CLK _25069_/D HRESETn VGND VGND VPWR VPWR _20739_/A sky130_fd_sc_hd__dfrtp_4
X_12034_ _11994_/Y _12019_/B _12019_/Y _12033_/X VGND VGND VPWR VPWR _12045_/A sky130_fd_sc_hd__a211o_4
X_16911_ _16940_/A VGND VGND VPWR VPWR _16936_/A sky130_fd_sc_hd__buf_2
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17891_ _17955_/A _17891_/B _17891_/C VGND VGND VPWR VPWR _17891_/X sky130_fd_sc_hd__and3_4
XFILLER_137_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19630_ _19628_/Y _19624_/X _19603_/X _19629_/X VGND VGND VPWR VPWR _19630_/X sky130_fd_sc_hd__a2bb2o_4
X_16842_ _16866_/A _16819_/Y _16841_/X VGND VGND VPWR VPWR _16852_/B sky130_fd_sc_hd__or3_4
XANTENNA__14087__B1 _13632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21028__D _21027_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19561_ _19559_/Y _19555_/X _11844_/X _19560_/X VGND VGND VPWR VPWR _23292_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13985_ _13971_/X _13984_/Y _13927_/A _13971_/X VGND VGND VPWR VPWR _24886_/D sky130_fd_sc_hd__a2bb2o_4
X_16773_ _16766_/X _16773_/B _16770_/X _16773_/D VGND VGND VPWR VPWR _16783_/C sky130_fd_sc_hd__or4_4
XFILLER_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18512_ _18486_/B _18507_/B _18475_/X _18509_/B VGND VGND VPWR VPWR _18513_/A sky130_fd_sc_hd__a211o_4
XFILLER_92_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12936_ _12854_/Y _12935_/X VGND VGND VPWR VPWR _12937_/A sky130_fd_sc_hd__or2_4
X_15724_ _15724_/A VGND VGND VPWR VPWR _24466_/D sky130_fd_sc_hd__inv_2
XFILLER_59_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15604__A _15604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19492_ _21939_/B _19489_/X _19445_/X _19489_/X VGND VGND VPWR VPWR _19492_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24566__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18443_ _18442_/A _18442_/B VGND VGND VPWR VPWR _18443_/Y sky130_fd_sc_hd__nand2_4
X_12867_ _12822_/X _12866_/X VGND VGND VPWR VPWR _12867_/X sky130_fd_sc_hd__or2_4
X_15655_ _15655_/A VGND VGND VPWR VPWR _22147_/A sky130_fd_sc_hd__buf_2
XANTENNA__15587__B1 _24532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11818_ _11818_/A VGND VGND VPWR VPWR _11818_/Y sky130_fd_sc_hd__inv_2
X_14606_ _23665_/D VGND VGND VPWR VPWR _20729_/B sky130_fd_sc_hd__inv_2
X_15586_ _15574_/X _15582_/X _15320_/X _24533_/Q _15585_/X VGND VGND VPWR VPWR _24533_/D
+ sky130_fd_sc_hd__a32o_4
X_18374_ _16450_/A _23822_/Q _16450_/Y _18532_/A VGND VGND VPWR VPWR _18374_/X sky130_fd_sc_hd__o22a_4
XFILLER_61_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12798_ _22605_/A _22595_/A _12796_/Y _12797_/Y VGND VGND VPWR VPWR _12808_/A sky130_fd_sc_hd__o22a_4
XFILLER_30_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _14444_/B _14521_/X _21376_/A _14536_/X VGND VGND VPWR VPWR _14537_/Y sky130_fd_sc_hd__a22oi_4
X_17325_ _17315_/Y _17325_/B _17325_/C VGND VGND VPWR VPWR _17348_/B sky130_fd_sc_hd__or3_4
X_11749_ _13232_/A VGND VGND VPWR VPWR _11749_/X sky130_fd_sc_hd__buf_2
XFILLER_105_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22872__A2 _22868_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14468_ _14493_/A VGND VGND VPWR VPWR _19862_/A sky130_fd_sc_hd__buf_2
X_17256_ _25214_/Q _24002_/Q _11550_/Y _17255_/Y VGND VGND VPWR VPWR _17259_/C sky130_fd_sc_hd__o22a_4
XFILLER_35_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13419_ _24928_/Q VGND VGND VPWR VPWR _13419_/Y sky130_fd_sc_hd__inv_2
X_16207_ _24293_/Q VGND VGND VPWR VPWR _16207_/Y sky130_fd_sc_hd__inv_2
X_17187_ _17187_/A VGND VGND VPWR VPWR _17187_/X sky130_fd_sc_hd__buf_2
X_14399_ _14390_/D VGND VGND VPWR VPWR _14399_/X sky130_fd_sc_hd__buf_2
X_16138_ _16138_/A VGND VGND VPWR VPWR _16138_/X sky130_fd_sc_hd__buf_2
XANTENNA__22172__A _12328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16069_ _16068_/Y _16064_/X _15765_/X _16064_/X VGND VGND VPWR VPWR _16069_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16170__A _16165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22900__A _22900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19828_ _19828_/A VGND VGND VPWR VPWR _19828_/X sky130_fd_sc_hd__buf_2
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14832__A2_N _14801_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19759_ _19759_/A VGND VGND VPWR VPWR _19759_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22770_ _12415_/A _22606_/X _17089_/A _22652_/X VGND VGND VPWR VPWR _22773_/B sky130_fd_sc_hd__a2bb2o_4
X_21721_ _22226_/A _21720_/X _14801_/Y _20757_/X VGND VGND VPWR VPWR _21721_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14847__A2_N _24137_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24236__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24440_ _24459_/CLK _24440_/D HRESETn VGND VGND VPWR VPWR _24440_/Q sky130_fd_sc_hd__dfrtp_4
X_21652_ _22745_/B _21641_/X _21642_/X _21651_/X VGND VGND VPWR VPWR _21653_/C sky130_fd_sc_hd__a211o_4
XANTENNA_clkbuf_5_10_0_HCLK_A clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20032__A2_N _20027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14250__B1 _14228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20603_ _20602_/X VGND VGND VPWR VPWR _20603_/X sky130_fd_sc_hd__buf_2
XANTENNA__21251__A _21251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16990__D _16989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24371_ _24385_/CLK _24371_/D HRESETn VGND VGND VPWR VPWR _22294_/A sky130_fd_sc_hd__dfrtp_4
X_21583_ _13324_/X _21582_/X VGND VGND VPWR VPWR _21583_/X sky130_fd_sc_hd__or2_4
X_23322_ _24750_/CLK _23322_/D VGND VGND VPWR VPWR _19477_/A sky130_fd_sc_hd__dfxtp_4
X_20534_ _20534_/A VGND VGND VPWR VPWR _20534_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20874__B2 _21093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23253_ _23278_/CLK _23253_/D VGND VGND VPWR VPWR _23253_/Q sky130_fd_sc_hd__dfxtp_4
X_20465_ _20465_/A VGND VGND VPWR VPWR _20465_/X sky130_fd_sc_hd__buf_2
XANTENNA__18560__A _18484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22204_ _12345_/X _22178_/X _16986_/A _22167_/A VGND VGND VPWR VPWR _22205_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16999__B _16996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23871__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23184_ _25050_/CLK _23184_/D VGND VGND VPWR VPWR _23184_/Q sky130_fd_sc_hd__dfxtp_4
X_20396_ _20396_/A _20393_/X _20396_/C VGND VGND VPWR VPWR _20396_/X sky130_fd_sc_hd__and3_4
XFILLER_134_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25095__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23800__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22135_ _17595_/C _22637_/A _24034_/Q _22121_/X VGND VGND VPWR VPWR _22136_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15502__B1 _24558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25024__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22066_ _14523_/A _22066_/B _22065_/X VGND VGND VPWR VPWR _22066_/X sky130_fd_sc_hd__or3_4
XFILLER_59_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21017_ _14486_/X _21016_/X _24746_/Q VGND VGND VPWR VPWR _21017_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_101_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13209__A _13136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13770_ _13770_/A _13770_/B _13716_/D _13778_/A VGND VGND VPWR VPWR _13771_/A sky130_fd_sc_hd__or4_4
X_22968_ _22968_/A _22968_/B VGND VGND VPWR VPWR _22978_/B sky130_fd_sc_hd__and2_4
XFILLER_15_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18755__B1 _18685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12721_ _12709_/B VGND VGND VPWR VPWR _12722_/B sky130_fd_sc_hd__inv_2
X_21919_ _21924_/A _19536_/Y VGND VGND VPWR VPWR _21919_/X sky130_fd_sc_hd__or2_4
X_24707_ _24671_/CLK _15009_/X HRESETn VGND VGND VPWR VPWR _24707_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22899_ _22637_/X _22896_/Y _22677_/A _22898_/X VGND VGND VPWR VPWR _22899_/X sky130_fd_sc_hd__a2bb2o_4
X_15440_ _15440_/A VGND VGND VPWR VPWR _15441_/B sky130_fd_sc_hd__inv_2
X_12652_ _12652_/A _12652_/B _12651_/X VGND VGND VPWR VPWR _12653_/C sky130_fd_sc_hd__or3_4
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24638_ _23762_/CLK _15264_/X HRESETn VGND VGND VPWR VPWR _13730_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22257__A _21051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _25199_/Q VGND VGND VPWR VPWR _11603_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15371_ _15371_/A VGND VGND VPWR VPWR _22408_/A sky130_fd_sc_hd__inv_2
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ _12581_/A _12582_/A _12581_/Y _12582_/Y VGND VGND VPWR VPWR _12583_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14792__B2 _24096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24569_ _24573_/CLK _15481_/X HRESETn VGND VGND VPWR VPWR _24569_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19180__B1 _19089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14322_ _14317_/B VGND VGND VPWR VPWR _14322_/Y sky130_fd_sc_hd__inv_2
X_17110_ _17101_/A _17104_/X _17109_/Y VGND VGND VPWR VPWR _24045_/D sky130_fd_sc_hd__and3_4
XFILLER_12_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11534_ _15916_/A VGND VGND VPWR VPWR _15920_/A sky130_fd_sc_hd__inv_2
X_18090_ _18089_/Y _11767_/X _18089_/A _17226_/X VGND VGND VPWR VPWR _18104_/A sky130_fd_sc_hd__o22a_4
XANTENNA__23959__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17041_ _17041_/A VGND VGND VPWR VPWR _17042_/D sky130_fd_sc_hd__inv_2
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ _14248_/Y VGND VGND VPWR VPWR _14253_/X sky130_fd_sc_hd__buf_2
XANTENNA__12933__D _12933_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13204_ _13204_/A _23602_/Q VGND VGND VPWR VPWR _13204_/X sky130_fd_sc_hd__or2_4
X_14184_ _24828_/Q _14171_/X _24827_/Q _14176_/X VGND VGND VPWR VPWR _14184_/X sky130_fd_sc_hd__o22a_4
XFILLER_87_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13135_ _13076_/A VGND VGND VPWR VPWR _13136_/A sky130_fd_sc_hd__buf_2
X_18992_ _22061_/B _18991_/X _15541_/X _18991_/X VGND VGND VPWR VPWR _23494_/D sky130_fd_sc_hd__a2bb2o_4
X_13066_ _23890_/Q VGND VGND VPWR VPWR _13076_/A sky130_fd_sc_hd__buf_2
X_17943_ _17732_/A _17943_/B _17942_/X VGND VGND VPWR VPWR _17943_/X sky130_fd_sc_hd__and3_4
XANTENNA__15318__B _20926_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_116_0_HCLK clkbuf_7_58_0_HCLK/X VGND VGND VPWR VPWR _24728_/CLK sky130_fd_sc_hd__clkbuf_1
X_12017_ _12016_/X VGND VGND VPWR VPWR _12017_/Y sky130_fd_sc_hd__inv_2
X_17874_ _17689_/X _17874_/B _17873_/X VGND VGND VPWR VPWR _17874_/X sky130_fd_sc_hd__and3_4
XFILLER_26_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_179_0_HCLK clkbuf_7_89_0_HCLK/X VGND VGND VPWR VPWR _24566_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21593__A2 _22840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22790__A1 _20819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19613_ _19613_/A VGND VGND VPWR VPWR _19613_/X sky130_fd_sc_hd__buf_2
XANTENNA__22790__B2 _22789_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24747__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16825_ _16825_/A VGND VGND VPWR VPWR _16825_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21336__A _21336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19544_ _21462_/B _19539_/X _11853_/X _19539_/X VGND VGND VPWR VPWR _23298_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16756_ _16756_/A _16756_/B _16756_/C _16756_/D VGND VGND VPWR VPWR _16756_/X sky130_fd_sc_hd__or4_4
XFILLER_19_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13968_ _23647_/D _13967_/Y _14257_/A _23647_/D VGND VGND VPWR VPWR _24891_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15707_ _15693_/X _15689_/X _15706_/X _24470_/Q _15661_/A VGND VGND VPWR VPWR _15707_/X
+ sky130_fd_sc_hd__a32o_4
X_12919_ _22826_/A _12919_/B VGND VGND VPWR VPWR _12921_/B sky130_fd_sc_hd__or2_4
X_19475_ _23323_/Q VGND VGND VPWR VPWR _19475_/Y sky130_fd_sc_hd__inv_2
X_13899_ _13862_/Y _13899_/B VGND VGND VPWR VPWR _13900_/B sky130_fd_sc_hd__nor2_4
X_16687_ _15938_/Y _17482_/A _15938_/Y _17482_/A VGND VGND VPWR VPWR _16687_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18426_ _18373_/A _18361_/A _18426_/C _18426_/D VGND VGND VPWR VPWR _18426_/X sky130_fd_sc_hd__or4_4
X_15638_ _15637_/X VGND VGND VPWR VPWR _21088_/A sky130_fd_sc_hd__inv_2
XFILLER_76_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22167__A _22167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18357_ _18357_/A _18357_/B _18357_/C _18356_/X VGND VGND VPWR VPWR _18378_/B sky130_fd_sc_hd__or4_4
X_15569_ _20806_/A VGND VGND VPWR VPWR _21292_/A sky130_fd_sc_hd__buf_2
XANTENNA__15980__B1 _15978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16165__A _16165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19171__B1 _19170_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12794__B1 _12793_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17308_ _17349_/A _17288_/Y VGND VGND VPWR VPWR _17308_/X sky130_fd_sc_hd__or2_4
XFILLER_30_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18288_ _18205_/D _18272_/B _18237_/X _18286_/B VGND VGND VPWR VPWR _18289_/A sky130_fd_sc_hd__a211o_4
XANTENNA__23629__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17239_ _17239_/A VGND VGND VPWR VPWR _17317_/D sky130_fd_sc_hd__inv_2
X_20250_ _20191_/B _20249_/X _20234_/X VGND VGND VPWR VPWR _20252_/C sky130_fd_sc_hd__o21a_4
XFILLER_116_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16288__A1 _15915_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20181_ _20193_/A _20192_/A _20158_/Y VGND VGND VPWR VPWR _20181_/X sky130_fd_sc_hd__and3_4
XFILLER_118_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_12_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_12_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_75_0_HCLK clkbuf_7_74_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_75_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__23022__A2 _15919_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23940_ _23343_/CLK _23940_/D HRESETn VGND VGND VPWR VPWR _23940_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18985__B1 _18938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24488__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21246__A _21245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23871_ _23859_/CLK _18249_/Y HRESETn VGND VGND VPWR VPWR _23871_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24417__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22822_ _22821_/X VGND VGND VPWR VPWR _22822_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18737__B1 _17199_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14786__A2_N _24096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22261__A1_N _12406_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22753_ _22753_/A _22587_/B VGND VGND VPWR VPWR _22753_/X sky130_fd_sc_hd__and2_4
XFILLER_20_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24070__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21704_ _21564_/A _21693_/X _20837_/X _21703_/X VGND VGND VPWR VPWR _21705_/C sky130_fd_sc_hd__a211o_4
X_22684_ _22539_/X _22682_/X _20777_/X _22683_/X VGND VGND VPWR VPWR _22685_/A sky130_fd_sc_hd__o22a_4
XFILLER_129_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24423_ _24620_/CLK _15838_/X HRESETn VGND VGND VPWR VPWR _24423_/Q sky130_fd_sc_hd__dfrtp_4
X_21635_ _17636_/A _21627_/X _21634_/X VGND VGND VPWR VPWR _21635_/X sky130_fd_sc_hd__or3_4
XANTENNA__15971__B1 _11594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16075__A _16075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24354_ _24333_/CLK _16049_/X HRESETn VGND VGND VPWR VPWR _16048_/A sky130_fd_sc_hd__dfrtp_4
X_21566_ _21566_/A _20818_/X VGND VGND VPWR VPWR _21569_/B sky130_fd_sc_hd__or2_4
XFILLER_138_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22805__A _22879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23305_ _23303_/CLK _19524_/X VGND VGND VPWR VPWR _23305_/Q sky130_fd_sc_hd__dfxtp_4
X_20517_ _20517_/A _13510_/B VGND VGND VPWR VPWR _20517_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__19386__A _19372_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24285_ _24138_/CLK _24285_/D HRESETn VGND VGND VPWR VPWR _24285_/Q sky130_fd_sc_hd__dfrtp_4
X_21497_ _21489_/Y _21496_/X _21192_/X VGND VGND VPWR VPWR _21538_/C sky130_fd_sc_hd__o21a_4
XANTENNA__12108__A _24574_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25205__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22524__B _22524_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23236_ _23292_/CLK _19719_/X VGND VGND VPWR VPWR _19716_/A sky130_fd_sc_hd__dfxtp_4
X_20448_ _13506_/A _13506_/B VGND VGND VPWR VPWR _20448_/X sky130_fd_sc_hd__or2_4
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11947__A _15414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23167_ _25106_/CLK _19902_/X VGND VGND VPWR VPWR _19901_/A sky130_fd_sc_hd__dfxtp_4
X_20379_ _15288_/Y _20367_/X _20358_/X _20378_/X VGND VGND VPWR VPWR _20380_/A sky130_fd_sc_hd__a211o_4
X_22118_ _22198_/A VGND VGND VPWR VPWR _22118_/X sky130_fd_sc_hd__buf_2
XFILLER_121_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23098_ _23258_/CLK _23098_/D VGND VGND VPWR VPWR _23098_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22221__B1 _21246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14940_ _14939_/Y _24267_/Q _14939_/Y _24267_/Q VGND VGND VPWR VPWR _14943_/C sky130_fd_sc_hd__a2bb2o_4
X_22049_ _21490_/X _13624_/Y _22048_/X VGND VGND VPWR VPWR _22049_/X sky130_fd_sc_hd__and3_4
XFILLER_125_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24840__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22772__B2 _22657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14871_ _14839_/Y _14844_/A VGND VGND VPWR VPWR _14871_/X sky130_fd_sc_hd__or2_4
XANTENNA__24158__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16610_ _16575_/A VGND VGND VPWR VPWR _16610_/X sky130_fd_sc_hd__buf_2
X_13822_ _13813_/Y _13822_/B VGND VGND VPWR VPWR _13822_/X sky130_fd_sc_hd__and2_4
XFILLER_29_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17590_ _17590_/A VGND VGND VPWR VPWR _17591_/B sky130_fd_sc_hd__inv_2
X_13753_ _13753_/A _13776_/C _13753_/C _13761_/B VGND VGND VPWR VPWR _13769_/C sky130_fd_sc_hd__or4_4
X_16541_ _16541_/A VGND VGND VPWR VPWR _21729_/A sky130_fd_sc_hd__inv_2
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12704_ _12704_/A _12704_/B VGND VGND VPWR VPWR _12705_/C sky130_fd_sc_hd__or2_4
X_19260_ _19260_/A VGND VGND VPWR VPWR _19260_/X sky130_fd_sc_hd__buf_2
XFILLER_108_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13684_ _13677_/X VGND VGND VPWR VPWR _13684_/Y sky130_fd_sc_hd__inv_2
X_16472_ _16471_/Y _16395_/X _16216_/X _16395_/X VGND VGND VPWR VPWR _16472_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14214__B1 _14213_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18211_ _18211_/A VGND VGND VPWR VPWR _18300_/A sky130_fd_sc_hd__inv_2
X_12635_ _12915_/C VGND VGND VPWR VPWR _12963_/A sky130_fd_sc_hd__buf_2
X_15423_ _15421_/X _15415_/Y _15416_/X _20550_/A _15422_/X VGND VGND VPWR VPWR _15423_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19191_ _19196_/A VGND VGND VPWR VPWR _19191_/X sky130_fd_sc_hd__buf_2
XANTENNA__15962__B1 _11576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15354_ _15352_/Y _15353_/X _11563_/X _15353_/X VGND VGND VPWR VPWR _15354_/X sky130_fd_sc_hd__a2bb2o_4
X_18142_ _18244_/A VGND VGND VPWR VPWR _18221_/A sky130_fd_sc_hd__inv_2
XFILLER_19_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23793__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ _24521_/Q VGND VGND VPWR VPWR _12566_/Y sky130_fd_sc_hd__inv_2
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11517_ _16475_/A _15916_/A VGND VGND VPWR VPWR _11537_/A sky130_fd_sc_hd__or2_4
X_14305_ _14302_/Y _14300_/X _14304_/X _14300_/X VGND VGND VPWR VPWR _24785_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23722__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15285_ _15285_/A VGND VGND VPWR VPWR _15285_/X sky130_fd_sc_hd__buf_2
X_18073_ _11729_/X _17230_/X _18072_/X _18065_/B VGND VGND VPWR VPWR _18073_/X sky130_fd_sc_hd__o22a_4
X_12497_ _12497_/A _12497_/B VGND VGND VPWR VPWR _12499_/B sky130_fd_sc_hd__or2_4
XANTENNA__22434__B _20749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14236_ _16376_/A VGND VGND VPWR VPWR _14236_/X sky130_fd_sc_hd__buf_2
X_17024_ _17089_/A VGND VGND VPWR VPWR _17077_/A sky130_fd_sc_hd__inv_2
XFILLER_116_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24999__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14167_ _14160_/A _14170_/B _14166_/Y VGND VGND VPWR VPWR _24834_/D sky130_fd_sc_hd__o21a_4
XFILLER_113_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13118_ _11732_/A VGND VGND VPWR VPWR _13122_/A sky130_fd_sc_hd__buf_2
XANTENNA__24928__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14098_ _14072_/A VGND VGND VPWR VPWR _14099_/A sky130_fd_sc_hd__inv_2
X_18975_ _18982_/A VGND VGND VPWR VPWR _18975_/X sky130_fd_sc_hd__buf_2
XANTENNA__22450__A _22450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20889__B _20759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13049_ _13049_/A _23206_/Q VGND VGND VPWR VPWR _13050_/C sky130_fd_sc_hd__or2_4
X_17926_ _17783_/A _17924_/X _17926_/C VGND VGND VPWR VPWR _17930_/B sky130_fd_sc_hd__and3_4
XFILLER_79_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24581__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17857_ _17889_/A _17857_/B _17857_/C VGND VGND VPWR VPWR _17857_/X sky130_fd_sc_hd__and3_4
XFILLER_113_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24510__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11592__A _25202_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16808_ _15892_/Y _24065_/Q _15902_/Y _24062_/Q VGND VGND VPWR VPWR _16808_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17788_ _17861_/A _23564_/Q VGND VGND VPWR VPWR _17788_/X sky130_fd_sc_hd__or2_4
X_19527_ _23303_/Q VGND VGND VPWR VPWR _19527_/Y sky130_fd_sc_hd__inv_2
X_16739_ _16739_/A _16739_/B _16739_/C _16739_/D VGND VGND VPWR VPWR _16739_/X sky130_fd_sc_hd__or4_4
X_19458_ _19440_/Y VGND VGND VPWR VPWR _19458_/X sky130_fd_sc_hd__buf_2
XANTENNA__14205__B1 _13665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18409_ _18448_/A VGND VGND VPWR VPWR _18484_/A sky130_fd_sc_hd__buf_2
X_19389_ _19389_/A VGND VGND VPWR VPWR _19389_/Y sky130_fd_sc_hd__inv_2
X_21420_ _24327_/Q _22154_/B _22351_/A VGND VGND VPWR VPWR _21420_/X sky130_fd_sc_hd__o21a_4
XANTENNA__13312__A _13092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13443__A1_N _13441_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21351_ _21169_/A _19250_/Y VGND VGND VPWR VPWR _21353_/B sky130_fd_sc_hd__or2_4
XFILLER_124_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15705__B1 _21567_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22344__B _16393_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20302_ _18622_/X VGND VGND VPWR VPWR _20315_/C sky130_fd_sc_hd__buf_2
X_24070_ _24623_/CLK _24070_/D HRESETn VGND VGND VPWR VPWR _16833_/A sky130_fd_sc_hd__dfrtp_4
X_21282_ _13525_/Y _21280_/X _13498_/Y _21562_/A VGND VGND VPWR VPWR _21282_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20057__A2 _15410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23021_ _24355_/Q _22859_/X _22864_/X VGND VGND VPWR VPWR _23021_/X sky130_fd_sc_hd__o21a_4
X_20233_ _20257_/B _20232_/X VGND VGND VPWR VPWR _20233_/X sky130_fd_sc_hd__or2_4
XFILLER_104_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24669__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20164_ _20164_/A _20164_/B _20162_/X _20163_/X VGND VGND VPWR VPWR _20165_/A sky130_fd_sc_hd__or4_4
XANTENNA__22360__A _21642_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16681__A1 _20919_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16681__B2 _16680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20095_ _23093_/Q VGND VGND VPWR VPWR _22106_/B sky130_fd_sc_hd__inv_2
X_24972_ _25186_/CLK _13479_/X HRESETn VGND VGND VPWR VPWR _13402_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22754__A1 _21561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22510__D _21033_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23923_ _23925_/CLK _23923_/D HRESETn VGND VGND VPWR VPWR _23923_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_44_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21407__C _21366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_162_0_HCLK clkbuf_7_81_0_HCLK/X VGND VGND VPWR VPWR _23156_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24251__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_5_0_HCLK clkbuf_7_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_23854_ _23845_/CLK _23854_/D HRESETn VGND VGND VPWR VPWR _23854_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_19_0_HCLK clkbuf_7_9_0_HCLK/X VGND VGND VPWR VPWR _24962_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22506__A1 _24340_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22805_ _22879_/A _22805_/B _22805_/C VGND VGND VPWR VPWR _22832_/A sky130_fd_sc_hd__and3_4
X_23785_ _23789_/CLK _23785_/D HRESETn VGND VGND VPWR VPWR _23785_/Q sky130_fd_sc_hd__dfrtp_4
X_20997_ _20991_/X _20996_/X _14485_/Y VGND VGND VPWR VPWR _20997_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_129_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22736_ _22736_/A _22957_/B VGND VGND VPWR VPWR _22736_/X sky130_fd_sc_hd__and2_4
XANTENNA__16197__B1 _15978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15944__B1 _11555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22667_ _16423_/Y _22551_/A _14779_/Y _22225_/A VGND VGND VPWR VPWR _22667_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19135__B1 _19089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12420_ _25101_/Q _12419_/Y VGND VGND VPWR VPWR _12422_/B sky130_fd_sc_hd__or2_4
X_24406_ _24590_/CLK _24406_/D HRESETn VGND VGND VPWR VPWR _24406_/Q sky130_fd_sc_hd__dfrtp_4
X_21618_ _18043_/A _21615_/X _21617_/X VGND VGND VPWR VPWR _21618_/X sky130_fd_sc_hd__and3_4
X_22598_ _22598_/A _21984_/X VGND VGND VPWR VPWR _22598_/X sky130_fd_sc_hd__or2_4
X_12351_ _12340_/X _12351_/B _12351_/C _12350_/X VGND VGND VPWR VPWR _12352_/D sky130_fd_sc_hd__or4_4
XFILLER_51_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21493__A1 _22018_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24337_ _24201_/CLK _24337_/D HRESETn VGND VGND VPWR VPWR _24337_/Q sky130_fd_sc_hd__dfrtp_4
X_21549_ _21549_/A _16042_/A VGND VGND VPWR VPWR _21549_/X sky130_fd_sc_hd__and2_4
X_15070_ _15067_/C _15079_/B VGND VGND VPWR VPWR _15071_/B sky130_fd_sc_hd__or2_4
X_12282_ _12261_/A _12282_/B _12281_/Y VGND VGND VPWR VPWR _25109_/D sky130_fd_sc_hd__and3_4
X_24268_ _24140_/CLK _16274_/X HRESETn VGND VGND VPWR VPWR _22399_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15711__A3 _15635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14021_ _16301_/A _20852_/A VGND VGND VPWR VPWR _14046_/A sky130_fd_sc_hd__or2_4
X_23219_ _23292_/CLK _19768_/X VGND VGND VPWR VPWR _19767_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_106_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24199_ _24197_/CLK _24199_/D HRESETn VGND VGND VPWR VPWR _16450_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21796__A2 _21113_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22270__A _22263_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24339__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13892__A _13908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18760_ _18760_/A VGND VGND VPWR VPWR _19100_/A sky130_fd_sc_hd__buf_2
X_15972_ _22294_/A VGND VGND VPWR VPWR _15972_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17711_ _17717_/A VGND VGND VPWR VPWR _17916_/A sky130_fd_sc_hd__buf_2
X_14923_ _24264_/Q VGND VGND VPWR VPWR _14923_/Y sky130_fd_sc_hd__inv_2
X_18691_ _18690_/X VGND VGND VPWR VPWR _18697_/A sky130_fd_sc_hd__inv_2
XFILLER_91_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17642_ _23939_/Q VGND VGND VPWR VPWR _17642_/Y sky130_fd_sc_hd__inv_2
X_14854_ _14712_/X _14833_/Y _14997_/A _14823_/Y VGND VGND VPWR VPWR _14855_/D sky130_fd_sc_hd__a2bb2o_4
X_13805_ _13845_/A VGND VGND VPWR VPWR _13811_/A sky130_fd_sc_hd__inv_2
X_17573_ _17497_/A _17570_/X VGND VGND VPWR VPWR _17573_/X sky130_fd_sc_hd__or2_4
X_11997_ _25144_/Q VGND VGND VPWR VPWR _11997_/Y sky130_fd_sc_hd__inv_2
X_14785_ _14785_/A VGND VGND VPWR VPWR _14870_/A sky130_fd_sc_hd__inv_2
XANTENNA__18195__A _18459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16708__A _23961_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19312_ _19304_/Y VGND VGND VPWR VPWR _19312_/X sky130_fd_sc_hd__buf_2
XANTENNA__22429__B _22429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16524_ _16522_/Y _16518_/X _16093_/X _16523_/X VGND VGND VPWR VPWR _24171_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15612__A _15585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23974__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13736_ _24640_/Q _13728_/A _13730_/A _24637_/Q VGND VGND VPWR VPWR _13737_/A sky130_fd_sc_hd__or4_4
XFILLER_72_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25198__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19243_ _19243_/A VGND VGND VPWR VPWR _21826_/B sky130_fd_sc_hd__inv_2
XANTENNA__23903__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16455_ HWDATA[8] VGND VGND VPWR VPWR _16455_/X sky130_fd_sc_hd__buf_2
XFILLER_31_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13667_ _13647_/Y VGND VGND VPWR VPWR _13667_/X sky130_fd_sc_hd__buf_2
XANTENNA__25127__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14228__A _16369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15406_ _15405_/Y _15401_/X _15291_/X _15401_/X VGND VGND VPWR VPWR _15406_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12618_ _12679_/C _24528_/Q _25057_/Q _12617_/Y VGND VGND VPWR VPWR _12622_/C sky130_fd_sc_hd__a2bb2o_4
X_19174_ _19174_/A VGND VGND VPWR VPWR _19174_/Y sky130_fd_sc_hd__inv_2
X_13598_ _13557_/A _13557_/B VGND VGND VPWR VPWR _13598_/Y sky130_fd_sc_hd__nand2_4
X_16386_ _16385_/Y _16308_/A _16216_/X _16308_/A VGND VGND VPWR VPWR _16386_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18125_ _18118_/A VGND VGND VPWR VPWR _18125_/X sky130_fd_sc_hd__buf_2
XFILLER_34_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12549_ _25062_/Q VGND VGND VPWR VPWR _12549_/Y sky130_fd_sc_hd__inv_2
X_15337_ _24610_/Q VGND VGND VPWR VPWR _15337_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12971__A _12933_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22164__B _22952_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18056_ _17446_/X _18061_/B _18055_/Y _21363_/A _17462_/Y VGND VGND VPWR VPWR _18056_/X
+ sky130_fd_sc_hd__a32o_4
X_15268_ _13742_/C _15250_/A _15240_/A _13754_/A _15251_/B VGND VGND VPWR VPWR _15268_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16360__B1 _16100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21362__A1_N _21357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17007_ _16207_/Y _17027_/A _24317_/Q _17022_/B VGND VGND VPWR VPWR _17007_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11587__A _11587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14219_ _20701_/A _14212_/X _14218_/X _14201_/X VGND VGND VPWR VPWR _24817_/D sky130_fd_sc_hd__a2bb2o_4
X_15199_ _14969_/Y _15219_/A VGND VGND VPWR VPWR _15216_/A sky130_fd_sc_hd__or2_4
XANTENNA__22984__A1 _24285_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24762__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14123__C1 _14122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18958_ _18958_/A VGND VGND VPWR VPWR _18958_/X sky130_fd_sc_hd__buf_2
XFILLER_119_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14674__B1 _14055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24009__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17909_ _17877_/A _23448_/Q VGND VGND VPWR VPWR _17909_/X sky130_fd_sc_hd__or2_4
XFILLER_39_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18889_ _18888_/Y _18884_/X _18795_/X _18884_/X VGND VGND VPWR VPWR _23530_/D sky130_fd_sc_hd__a2bb2o_4
X_20920_ _20910_/X _20916_/X _20918_/X _20919_/X VGND VGND VPWR VPWR _20920_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_235_0_HCLK clkbuf_8_235_0_HCLK/A VGND VGND VPWR VPWR _23716_/CLK sky130_fd_sc_hd__clkbuf_1
X_20851_ _17219_/Y _17222_/B _21079_/B _20850_/Y VGND VGND VPWR VPWR _20852_/B sky130_fd_sc_hd__o22a_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16752__A2_N _16846_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15522__A _11630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23570_ _23560_/CLK _23570_/D VGND VGND VPWR VPWR _17860_/B sky130_fd_sc_hd__dfxtp_4
X_20782_ _20782_/A VGND VGND VPWR VPWR _20782_/X sky130_fd_sc_hd__buf_2
XPHY_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22521_ _22521_/A _21984_/X VGND VGND VPWR VPWR _22521_/X sky130_fd_sc_hd__or2_4
XANTENNA__23644__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15926__B1 _11522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22452_ _20926_/A VGND VGND VPWR VPWR _22452_/X sky130_fd_sc_hd__buf_2
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21403_ _21403_/A _21402_/X VGND VGND VPWR VPWR _21403_/X sky130_fd_sc_hd__and2_4
X_25171_ _23112_/CLK _25171_/D HRESETn VGND VGND VPWR VPWR _11850_/A sky130_fd_sc_hd__dfrtp_4
X_22383_ _20909_/X _22382_/X _22240_/X _11587_/A _21402_/X VGND VGND VPWR VPWR _22383_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_136_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24122_ _24113_/CLK _16630_/X HRESETn VGND VGND VPWR VPWR _14740_/A sky130_fd_sc_hd__dfrtp_4
X_21334_ _21144_/A _21334_/B _21334_/C VGND VGND VPWR VPWR _21334_/X sky130_fd_sc_hd__and3_4
XANTENNA__17168__B _16858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24053_ _24612_/CLK _17075_/Y HRESETn VGND VGND VPWR VPWR _24053_/Q sky130_fd_sc_hd__dfrtp_4
X_21265_ _20815_/X _21265_/B VGND VGND VPWR VPWR _21265_/X sky130_fd_sc_hd__and2_4
XFILLER_137_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22802__B _22745_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23004_ _23004_/A _23003_/X VGND VGND VPWR VPWR _23004_/X sky130_fd_sc_hd__and2_4
X_20216_ _20227_/A VGND VGND VPWR VPWR _20216_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16103__B1 _15788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21196_ _21238_/A VGND VGND VPWR VPWR _21367_/A sky130_fd_sc_hd__buf_2
XFILLER_46_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20603__A _20602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24432__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20147_ _20147_/A VGND VGND VPWR VPWR _20147_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_45_0_HCLK clkbuf_6_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_91_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20078_ _22084_/B _20077_/X _19597_/A _20077_/X VGND VGND VPWR VPWR _20078_/X sky130_fd_sc_hd__a2bb2o_4
X_24955_ _24824_/CLK _24955_/D HRESETn VGND VGND VPWR VPWR _11679_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11920_ _22030_/A _11919_/X _25163_/Q _11919_/X VGND VGND VPWR VPWR _25164_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23906_ _23908_/CLK _18014_/X HRESETn VGND VGND VPWR VPWR _23906_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12121__A _24562_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24886_ _23774_/CLK _24886_/D HRESETn VGND VGND VPWR VPWR _13927_/A sky130_fd_sc_hd__dfrtp_4
X_11851_ _19614_/A VGND VGND VPWR VPWR _11851_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21434__A _21434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14968__B2 _24259_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23837_ _23828_/CLK _23837_/D HRESETn VGND VGND VPWR VPWR _23837_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19356__B1 _19311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15432__A _15431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14570_ _17717_/A VGND VGND VPWR VPWR _17742_/A sky130_fd_sc_hd__buf_2
X_11782_ _11780_/Y _11828_/B _13551_/B VGND VGND VPWR VPWR _11782_/X sky130_fd_sc_hd__o21a_4
XFILLER_14_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23768_ _24728_/CLK _20243_/X HRESETn VGND VGND VPWR VPWR _20254_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__16709__A2 _23961_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_HCLK clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_13521_ _13521_/A VGND VGND VPWR VPWR _13521_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22719_ _11557_/Y _22536_/X _15945_/Y _22537_/X VGND VGND VPWR VPWR _22719_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25220__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23699_ _24162_/CLK _20436_/Y HRESETn VGND VGND VPWR VPWR _13503_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18743__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13452_ _24938_/Q _14387_/C _13450_/Y _14394_/A VGND VGND VPWR VPWR _13453_/D sky130_fd_sc_hd__o22a_4
X_16240_ _16240_/A VGND VGND VPWR VPWR _16256_/A sky130_fd_sc_hd__inv_2
XFILLER_9_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22265__A _14897_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12403_ _12508_/A _12403_/B VGND VGND VPWR VPWR _12409_/B sky130_fd_sc_hd__or2_4
XFILLER_40_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13383_ _11916_/X VGND VGND VPWR VPWR _20691_/B sky130_fd_sc_hd__buf_2
X_16171_ _16169_/Y _16165_/X _15772_/X _16170_/X VGND VGND VPWR VPWR _16171_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12334_ _25077_/Q VGND VGND VPWR VPWR _12407_/B sky130_fd_sc_hd__inv_2
X_15122_ _15154_/A _15120_/X _15121_/X VGND VGND VPWR VPWR _15122_/X sky130_fd_sc_hd__and3_4
XANTENNA__16342__B1 _16264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15053_ _15019_/A _15051_/A VGND VGND VPWR VPWR _15054_/C sky130_fd_sc_hd__or2_4
X_19930_ _21943_/B _19927_/X _19445_/A _19927_/X VGND VGND VPWR VPWR _23157_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_127_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_255_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12265_ _12265_/A _12265_/B _12265_/C _12298_/A VGND VGND VPWR VPWR _12265_/X sky130_fd_sc_hd__or4_4
XFILLER_120_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14004_ _24809_/Q VGND VGND VPWR VPWR _14004_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_6_0_HCLK_A clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19861_ _23182_/Q VGND VGND VPWR VPWR _22071_/B sky130_fd_sc_hd__inv_2
X_12196_ _12154_/Y _12193_/X _12188_/B _12195_/X VGND VGND VPWR VPWR _12196_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24173__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18812_ _18811_/Y _18809_/X _18740_/X _18809_/X VGND VGND VPWR VPWR _23557_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15607__A _15604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19792_ _19792_/A VGND VGND VPWR VPWR _19792_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24102__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18743_ HWDATA[5] VGND VGND VPWR VPWR _18743_/X sky130_fd_sc_hd__buf_2
X_15955_ _22598_/A VGND VGND VPWR VPWR _15955_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12667__C1 _12666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14906_ _24669_/Q VGND VGND VPWR VPWR _15105_/A sky130_fd_sc_hd__inv_2
XFILLER_3_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18674_ _18672_/Y _18668_/X _17205_/X _18673_/X VGND VGND VPWR VPWR _18674_/X sky130_fd_sc_hd__a2bb2o_4
X_15886_ _15884_/Y _15880_/X _15511_/X _15885_/X VGND VGND VPWR VPWR _24404_/D sky130_fd_sc_hd__a2bb2o_4
X_17625_ _17625_/A VGND VGND VPWR VPWR _17625_/Y sky130_fd_sc_hd__inv_2
X_14837_ _24686_/Q _14835_/Y _24688_/Q _14836_/Y VGND VGND VPWR VPWR _14837_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14959__B2 _14958_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15620__A2 _15617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17556_ _17497_/D _17550_/X _17520_/X _17553_/B VGND VGND VPWR VPWR _17556_/X sky130_fd_sc_hd__a211o_4
XFILLER_17_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_65_0_HCLK clkbuf_8_65_0_HCLK/A VGND VGND VPWR VPWR _24840_/CLK sky130_fd_sc_hd__clkbuf_1
X_14768_ _24699_/Q VGND VGND VPWR VPWR _15034_/A sky130_fd_sc_hd__inv_2
XFILLER_32_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16507_ _16505_/Y _16506_/X _16259_/X _16506_/X VGND VGND VPWR VPWR _24178_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13719_ _13718_/X VGND VGND VPWR VPWR _13780_/B sky130_fd_sc_hd__buf_2
X_17487_ _23945_/Q VGND VGND VPWR VPWR _17487_/Y sky130_fd_sc_hd__inv_2
X_14699_ _24099_/Q VGND VGND VPWR VPWR _14699_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19226_ _19212_/Y VGND VGND VPWR VPWR _19226_/X sky130_fd_sc_hd__buf_2
X_16438_ _16438_/A VGND VGND VPWR VPWR _16438_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13395__B1 SCLK_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19157_ _23434_/Q VGND VGND VPWR VPWR _19157_/Y sky130_fd_sc_hd__inv_2
X_16369_ _16369_/A VGND VGND VPWR VPWR _16369_/X sky130_fd_sc_hd__buf_2
XFILLER_8_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18108_ _18093_/A VGND VGND VPWR VPWR _18108_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24943__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19088_ _23458_/Q VGND VGND VPWR VPWR _19088_/Y sky130_fd_sc_hd__inv_2
X_18039_ _18038_/X VGND VGND VPWR VPWR _18039_/X sky130_fd_sc_hd__buf_2
X_21050_ _15576_/X VGND VGND VPWR VPWR _21050_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21519__A _21519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20001_ _20000_/Y _19996_/X _15522_/X _19996_/X VGND VGND VPWR VPWR _23130_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18828__A _18711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17732__A _17732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21952_ _21948_/X _21951_/X _14524_/D VGND VGND VPWR VPWR _21952_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_39_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23896__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24740_ _24740_/CLK _14550_/X HRESETn VGND VGND VPWR VPWR _24740_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12390__A2_N _24470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20903_ _20902_/X VGND VGND VPWR VPWR _20903_/X sky130_fd_sc_hd__buf_2
XANTENNA__16691__A2_N _17490_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23825__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24671_ _24671_/CLK _15165_/X HRESETn VGND VGND VPWR VPWR _24671_/Q sky130_fd_sc_hd__dfrtp_4
X_21883_ _16459_/Y _21882_/X _24099_/Q _21570_/A VGND VGND VPWR VPWR _21883_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15072__B1 _14984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25049__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23622_ _24783_/CLK _20714_/X HRESETn VGND VGND VPWR VPWR _23622_/Q sky130_fd_sc_hd__dfrtp_4
X_20834_ _20834_/A _22228_/A VGND VGND VPWR VPWR _20834_/Y sky130_fd_sc_hd__nor2_4
XFILLER_42_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23553_ _24998_/CLK _23553_/D VGND VGND VPWR VPWR _13226_/B sky130_fd_sc_hd__dfxtp_4
X_20765_ _21357_/A _20764_/X _18130_/Y _21357_/A VGND VGND VPWR VPWR _20765_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19659__A _19646_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22504_ _14812_/A _22147_/X _22148_/X _22503_/X VGND VGND VPWR VPWR _22504_/X sky130_fd_sc_hd__a211o_4
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23484_ _23486_/CLK _23484_/D VGND VGND VPWR VPWR _23484_/Q sky130_fd_sc_hd__dfxtp_4
X_20696_ _20696_/A _20697_/B VGND VGND VPWR VPWR _23796_/D sky130_fd_sc_hd__and2_4
XANTENNA__16572__B1 _16243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22435_ _20832_/A VGND VGND VPWR VPWR _22435_/X sky130_fd_sc_hd__buf_2
XFILLER_13_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24684__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25154_ _24953_/CLK _25154_/D HRESETn VGND VGND VPWR VPWR _25154_/Q sky130_fd_sc_hd__dfrtp_4
X_22366_ _22198_/A VGND VGND VPWR VPWR _22366_/X sky130_fd_sc_hd__buf_2
XANTENNA__16324__B1 _15479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24613__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24105_ _24112_/CLK _24105_/D HRESETn VGND VGND VPWR VPWR _24105_/Q sky130_fd_sc_hd__dfrtp_4
X_21317_ _24014_/Q _15653_/X _21314_/X _21315_/X _21316_/X VGND VGND VPWR VPWR _21318_/A
+ sky130_fd_sc_hd__a2111o_4
X_25085_ _25091_/CLK _25085_/D HRESETn VGND VGND VPWR VPWR _12373_/A sky130_fd_sc_hd__dfrtp_4
X_22297_ _24440_/Q _20787_/B VGND VGND VPWR VPWR _22297_/X sky130_fd_sc_hd__or2_4
XFILLER_117_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12050_ _12045_/X VGND VGND VPWR VPWR _20693_/B sky130_fd_sc_hd__inv_2
X_24036_ _24031_/CLK _24036_/D HRESETn VGND VGND VPWR VPWR _16986_/A sky130_fd_sc_hd__dfrtp_4
X_21248_ _13358_/X VGND VGND VPWR VPWR _21248_/X sky130_fd_sc_hd__buf_2
XFILLER_46_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12897__C1 _12896_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11955__A _16301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12361__B2 _22373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15427__A _15426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21179_ _21179_/A VGND VGND VPWR VPWR _21400_/A sky130_fd_sc_hd__buf_2
XFILLER_132_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23066__D _20413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24021__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15740_ _15740_/A VGND VGND VPWR VPWR _15740_/X sky130_fd_sc_hd__buf_2
X_12952_ _12952_/A _12947_/X _12952_/C VGND VGND VPWR VPWR _12952_/X sky130_fd_sc_hd__and3_4
X_24938_ _24968_/CLK _24938_/D HRESETn VGND VGND VPWR VPWR _24938_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11903_ _22006_/A _11886_/X _11887_/Y _11902_/X VGND VGND VPWR VPWR _11903_/X sky130_fd_sc_hd__a211o_4
X_15671_ _15658_/X _15647_/X _15477_/X _24493_/Q _15661_/X VGND VGND VPWR VPWR _24493_/D
+ sky130_fd_sc_hd__a32o_4
X_12883_ _12933_/D _12883_/B VGND VGND VPWR VPWR _12883_/X sky130_fd_sc_hd__or2_4
X_24869_ _23680_/CLK _24869_/D HRESETn VGND VGND VPWR VPWR _24869_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_73_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17410_ _17273_/Y _17429_/A VGND VGND VPWR VPWR _17411_/B sky130_fd_sc_hd__or2_4
X_14622_ _14620_/A VGND VGND VPWR VPWR _14622_/X sky130_fd_sc_hd__buf_2
X_11834_ _19600_/A VGND VGND VPWR VPWR _11834_/Y sky130_fd_sc_hd__inv_2
X_18390_ _16430_/Y _18503_/A _24211_/Q _18491_/A VGND VGND VPWR VPWR _18390_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14810__B1 _15003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17340_/X VGND VGND VPWR VPWR _17342_/B sky130_fd_sc_hd__inv_2
XFILLER_57_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18001__B1 _23913_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11765_ _11765_/A _11728_/X VGND VGND VPWR VPWR _11765_/X sky130_fd_sc_hd__or2_4
X_14553_ _19946_/B VGND VGND VPWR VPWR _14553_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _20438_/A _13503_/X VGND VGND VPWR VPWR _13505_/B sky130_fd_sc_hd__or2_4
XPHY_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17272_ _23979_/Q VGND VGND VPWR VPWR _17323_/C sky130_fd_sc_hd__inv_2
XFILLER_41_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _11708_/B _11718_/B VGND VGND VPWR VPWR _11696_/X sky130_fd_sc_hd__or2_4
X_14484_ _14479_/A VGND VGND VPWR VPWR _14484_/X sky130_fd_sc_hd__buf_2
XPHY_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19011_ _14540_/X _19862_/B _19509_/C VGND VGND VPWR VPWR _19012_/A sky130_fd_sc_hd__or3_4
XFILLER_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16223_ _16223_/A VGND VGND VPWR VPWR _16223_/Y sky130_fd_sc_hd__inv_2
X_13435_ _13435_/A VGND VGND VPWR VPWR _13435_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21439__B2 _13333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14506__A _14480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13366_ _13363_/A VGND VGND VPWR VPWR _13366_/X sky130_fd_sc_hd__buf_2
X_16154_ _16151_/Y _16152_/X _16153_/X _16152_/X VGND VGND VPWR VPWR _24315_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16315__B1 _16243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14225__B _18633_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24354__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15105_ _15105_/A _15179_/A _14950_/Y _14941_/Y VGND VGND VPWR VPWR _15105_/X sky130_fd_sc_hd__or4_4
X_12317_ _12317_/A VGND VGND VPWR VPWR _12416_/A sky130_fd_sc_hd__inv_2
X_13297_ _13297_/A _23069_/Q VGND VGND VPWR VPWR _13297_/X sky130_fd_sc_hd__or2_4
X_16085_ _16082_/Y _16084_/X _11576_/X _16084_/X VGND VGND VPWR VPWR _24340_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12248_ _12083_/X _12252_/B VGND VGND VPWR VPWR _12249_/C sky130_fd_sc_hd__nand2_4
X_15036_ _15018_/X _15036_/B _15035_/Y VGND VGND VPWR VPWR _24700_/D sky130_fd_sc_hd__and3_4
X_19913_ _23163_/Q VGND VGND VPWR VPWR _21677_/B sky130_fd_sc_hd__inv_2
XFILLER_138_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21339__A _21339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19844_ _23189_/Q VGND VGND VPWR VPWR _21950_/B sky130_fd_sc_hd__inv_2
XFILLER_9_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15337__A _24610_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12179_ _12299_/A VGND VGND VPWR VPWR _12265_/C sky130_fd_sc_hd__inv_2
XFILLER_111_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19775_ _19774_/Y _19772_/X _19731_/X _19772_/X VGND VGND VPWR VPWR _23216_/D sky130_fd_sc_hd__a2bb2o_4
X_16987_ _16195_/A _16986_/A _16195_/Y _17034_/A VGND VGND VPWR VPWR _16987_/X sky130_fd_sc_hd__o22a_4
XFILLER_111_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18726_ _17888_/B VGND VGND VPWR VPWR _18726_/Y sky130_fd_sc_hd__inv_2
X_15938_ _22820_/A VGND VGND VPWR VPWR _15938_/Y sky130_fd_sc_hd__inv_2
X_18657_ _18644_/Y VGND VGND VPWR VPWR _18657_/X sky130_fd_sc_hd__buf_2
X_15869_ _15866_/Y _15868_/X _11576_/X _15868_/X VGND VGND VPWR VPWR _15869_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25142__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17608_ _17587_/X VGND VGND VPWR VPWR _17609_/B sky130_fd_sc_hd__inv_2
X_18588_ _16328_/Y _18479_/A _16328_/Y _18479_/A VGND VGND VPWR VPWR _18592_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17539_ _16702_/Y _17534_/B _17520_/X _17535_/Y VGND VGND VPWR VPWR _17539_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22875__B1 _22874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20550_ _20550_/A VGND VGND VPWR VPWR _20554_/A sky130_fd_sc_hd__inv_2
XANTENNA__16554__B1 _16216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_9_0_HCLK clkbuf_6_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__20418__A _20425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19209_ _23415_/Q VGND VGND VPWR VPWR _19209_/Y sky130_fd_sc_hd__inv_2
X_20481_ _13509_/B _13509_/C VGND VGND VPWR VPWR _20481_/X sky130_fd_sc_hd__or2_4
X_22220_ _20457_/Y _20927_/X _20594_/Y _21870_/A VGND VGND VPWR VPWR _22220_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24095__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22151_ _11680_/Y _20940_/X _24933_/Q _13630_/C VGND VGND VPWR VPWR _22151_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17727__A _17727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21102_ _16621_/A _21095_/X _21099_/X _21100_/X _21101_/X VGND VGND VPWR VPWR _21103_/A
+ sky130_fd_sc_hd__a32o_4
X_22082_ _14471_/A _22074_/X _22082_/C VGND VGND VPWR VPWR _22082_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_110_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_221_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21033_ _11939_/A _15407_/Y _21088_/A _15424_/Y VGND VGND VPWR VPWR _21033_/X sky130_fd_sc_hd__or4_4
XFILLER_82_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18558__A _18484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22984_ _24285_/Q _22859_/X _22338_/A VGND VGND VPWR VPWR _22984_/X sky130_fd_sc_hd__o21a_4
X_24723_ _24723_/CLK _14663_/X HRESETn VGND VGND VPWR VPWR _24723_/Q sky130_fd_sc_hd__dfrtp_4
X_21935_ _21935_/A _21935_/B VGND VGND VPWR VPWR _21936_/C sky130_fd_sc_hd__or2_4
XFILLER_76_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16078__A _16078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21866_ _13532_/A VGND VGND VPWR VPWR _21866_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24654_ _24654_/CLK _24654_/D HRESETn VGND VGND VPWR VPWR _14955_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _22971_/A _20778_/X _20795_/X _20811_/X _20816_/X VGND VGND VPWR VPWR _21028_/B
+ sky130_fd_sc_hd__a32o_4
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23605_ _24005_/CLK _23605_/D VGND VGND VPWR VPWR _18670_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22866__B1 _21694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21797_ _21796_/X VGND VGND VPWR VPWR _21797_/Y sky130_fd_sc_hd__inv_2
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24585_ _24587_/CLK _15404_/X HRESETn VGND VGND VPWR VPWR _24585_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ _25214_/Q VGND VGND VPWR VPWR _11550_/Y sky130_fd_sc_hd__inv_2
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20748_ _20747_/X VGND VGND VPWR VPWR _20748_/X sky130_fd_sc_hd__buf_2
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23536_ _23537_/CLK _23536_/D VGND VGND VPWR VPWR _13259_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_23_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23467_ _23416_/CLK _19067_/X VGND VGND VPWR VPWR _17812_/B sky130_fd_sc_hd__dfxtp_4
X_20679_ _23757_/Q VGND VGND VPWR VPWR _20679_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13220_ _13110_/A _19477_/A VGND VGND VPWR VPWR _13221_/C sky130_fd_sc_hd__or2_4
XANTENNA__16560__A3 _16558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22418_ _22163_/A VGND VGND VPWR VPWR _22418_/X sky130_fd_sc_hd__buf_2
X_25206_ _24372_/CLK _25206_/D HRESETn VGND VGND VPWR VPWR _11575_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_137_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23398_ _25194_/CLK _19262_/X VGND VGND VPWR VPWR _22047_/A sky130_fd_sc_hd__dfxtp_4
X_13151_ _13026_/X _13147_/X _13151_/C VGND VGND VPWR VPWR _13151_/X sky130_fd_sc_hd__or3_4
XFILLER_87_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22349_ _16443_/A _22349_/B VGND VGND VPWR VPWR _22349_/X sky130_fd_sc_hd__or2_4
XFILLER_128_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25137_ _24840_/CLK _12052_/X HRESETn VGND VGND VPWR VPWR _25137_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20845__A2_N _14015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12102_ _25126_/Q _24569_/Q _12219_/A _12101_/Y VGND VGND VPWR VPWR _12106_/C sky130_fd_sc_hd__o22a_4
X_13082_ _13076_/A VGND VGND VPWR VPWR _13204_/A sky130_fd_sc_hd__buf_2
XANTENNA__23043__B1 _25221_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25068_ _25061_/CLK _25068_/D HRESETn VGND VGND VPWR VPWR _25068_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12033_ _12023_/X _12024_/X _12028_/X _12033_/D VGND VGND VPWR VPWR _12033_/X sky130_fd_sc_hd__or4_4
X_16910_ _16910_/A VGND VGND VPWR VPWR _24073_/D sky130_fd_sc_hd__inv_2
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24019_ _23676_/CLK _24019_/D HRESETn VGND VGND VPWR VPWR _20396_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_2_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17890_ _17738_/A _17890_/B _17889_/X VGND VGND VPWR VPWR _17891_/C sky130_fd_sc_hd__or3_4
XFILLER_132_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16841_ _16863_/A _16769_/Y _16822_/X _16841_/D VGND VGND VPWR VPWR _16841_/X sky130_fd_sc_hd__or4_4
XANTENNA__23747__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_15_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19560_ _19554_/Y VGND VGND VPWR VPWR _19560_/X sky130_fd_sc_hd__buf_2
XFILLER_120_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16772_ _15889_/A _16771_/A _15889_/Y _16771_/Y VGND VGND VPWR VPWR _16773_/D sky130_fd_sc_hd__o22a_4
X_13984_ _13956_/X _13983_/X _14230_/A _13963_/X VGND VGND VPWR VPWR _13984_/Y sky130_fd_sc_hd__a22oi_4
X_18511_ _18504_/A _18511_/B _18511_/C VGND VGND VPWR VPWR _23828_/D sky130_fd_sc_hd__and3_4
X_15723_ _15712_/X _15713_/X _13474_/B _15717_/C _15722_/X VGND VGND VPWR VPWR _15724_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_59_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12935_ _12881_/X _12943_/D VGND VGND VPWR VPWR _12935_/X sky130_fd_sc_hd__or2_4
X_19491_ _19491_/A VGND VGND VPWR VPWR _21939_/B sky130_fd_sc_hd__inv_2
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18442_ _18442_/A _18442_/B VGND VGND VPWR VPWR _18444_/B sky130_fd_sc_hd__or2_4
X_15654_ _15653_/X VGND VGND VPWR VPWR _15655_/A sky130_fd_sc_hd__buf_2
X_12866_ _12835_/X _12844_/X _12866_/C _12865_/X VGND VGND VPWR VPWR _12866_/X sky130_fd_sc_hd__or4_4
XFILLER_18_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14605_ _18759_/B _16035_/B _19167_/B VGND VGND VPWR VPWR _24731_/D sky130_fd_sc_hd__o21a_4
X_11817_ _11817_/A _11817_/B VGND VGND VPWR VPWR _11817_/X sky130_fd_sc_hd__and2_4
X_18373_ _18373_/A VGND VGND VPWR VPWR _18532_/A sky130_fd_sc_hd__buf_2
X_15585_ _15585_/A VGND VGND VPWR VPWR _15585_/X sky130_fd_sc_hd__buf_2
X_12797_ _22595_/A VGND VGND VPWR VPWR _12797_/Y sky130_fd_sc_hd__inv_2
XPHY_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17324_/A _17324_/B _17324_/C VGND VGND VPWR VPWR _17325_/C sky130_fd_sc_hd__or3_4
X_14536_ _21378_/A _14526_/Y VGND VGND VPWR VPWR _14536_/X sky130_fd_sc_hd__or2_4
XPHY_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _11733_/A VGND VGND VPWR VPWR _13232_/A sky130_fd_sc_hd__buf_2
XANTENNA__16536__B1 _16455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12963__B _12933_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24535__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_139_0_HCLK clkbuf_7_69_0_HCLK/X VGND VGND VPWR VPWR _23482_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17255_ _24002_/Q VGND VGND VPWR VPWR _17255_/Y sky130_fd_sc_hd__inv_2
X_14467_ _24742_/Q VGND VGND VPWR VPWR _14493_/A sky130_fd_sc_hd__buf_2
X_11679_ _11679_/A VGND VGND VPWR VPWR _11679_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14236__A _16376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16206_ _16205_/Y _16203_/X _15897_/X _16203_/X VGND VGND VPWR VPWR _16206_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13418_ _13418_/A _13418_/B _13414_/X _13418_/D VGND VGND VPWR VPWR _13454_/A sky130_fd_sc_hd__or4_4
X_17186_ _17186_/A _17186_/B VGND VGND VPWR VPWR _17187_/A sky130_fd_sc_hd__or2_4
X_14398_ _14393_/Y _14371_/X _14397_/X _13608_/X _14387_/A VGND VGND VPWR VPWR _14398_/X
+ sky130_fd_sc_hd__a32o_4
X_16137_ _16137_/A VGND VGND VPWR VPWR _16138_/A sky130_fd_sc_hd__buf_2
X_13349_ _13348_/Y _13344_/X _11631_/X _13344_/X VGND VGND VPWR VPWR _24990_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23647__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16451__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16068_ _24346_/Q VGND VGND VPWR VPWR _16068_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15019_ _15019_/A _15019_/B _14878_/A _14974_/X VGND VGND VPWR VPWR _15019_/X sky130_fd_sc_hd__or4_4
XANTENNA__21596__B1 _21113_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19827_ _23194_/Q VGND VGND VPWR VPWR _21525_/B sky130_fd_sc_hd__inv_2
XFILLER_111_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19758_ _19531_/A _18038_/X _19530_/A _19644_/X VGND VGND VPWR VPWR _19759_/A sky130_fd_sc_hd__or4_4
XFILLER_49_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18709_ _18708_/Y _18705_/X _18685_/X _18705_/X VGND VGND VPWR VPWR _23592_/D sky130_fd_sc_hd__a2bb2o_4
X_19689_ _19688_/Y VGND VGND VPWR VPWR _19689_/X sky130_fd_sc_hd__buf_2
XFILLER_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21720_ _14937_/Y _21720_/B VGND VGND VPWR VPWR _21720_/X sky130_fd_sc_hd__and2_4
XANTENNA__19961__B1 _19387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21651_ _15824_/A _21651_/B VGND VGND VPWR VPWR _21651_/X sky130_fd_sc_hd__and2_4
XANTENNA__16661__A1_N _14709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_35_0_HCLK clkbuf_7_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_71_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20602_ _20651_/A VGND VGND VPWR VPWR _20602_/X sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_4_9_0_HCLK_A clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21251__B _20826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24370_ _24385_/CLK _24370_/D HRESETn VGND VGND VPWR VPWR _22239_/A sky130_fd_sc_hd__dfrtp_4
X_21582_ _20847_/A _20758_/X VGND VGND VPWR VPWR _21582_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_98_0_HCLK clkbuf_7_99_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_98_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__21520__B1 _21231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24276__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23321_ _24750_/CLK _19481_/X VGND VGND VPWR VPWR _23321_/Q sky130_fd_sc_hd__dfxtp_4
X_20533_ _20511_/X _20532_/Y _24610_/Q _20515_/X VGND VGND VPWR VPWR _20533_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12375__A1_N _12489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24205__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23252_ _23242_/CLK _19674_/X VGND VGND VPWR VPWR _23252_/Q sky130_fd_sc_hd__dfxtp_4
X_20464_ _20414_/X VGND VGND VPWR VPWR _20465_/A sky130_fd_sc_hd__inv_2
XFILLER_14_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22363__A _22438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22203_ _22203_/A _22163_/A VGND VGND VPWR VPWR _22203_/X sky130_fd_sc_hd__and2_4
XFILLER_119_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20087__B1 _19610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23183_ _25050_/CLK _19860_/X VGND VGND VPWR VPWR _19858_/A sky130_fd_sc_hd__dfxtp_4
X_20395_ _23678_/Q _17182_/B _20394_/Y _20343_/Y VGND VGND VPWR VPWR _20396_/C sky130_fd_sc_hd__a211o_4
Xclkbuf_3_4_0_HCLK clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22134_ _25077_/Q _20814_/X VGND VGND VPWR VPWR _22136_/C sky130_fd_sc_hd__and2_4
XFILLER_82_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22065_ _21665_/A _22063_/X _22065_/C VGND VGND VPWR VPWR _22065_/X sky130_fd_sc_hd__and3_4
XFILLER_138_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22810__B _22884_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21016_ _14528_/A _21012_/X _21013_/X _21014_/X _21015_/X VGND VGND VPWR VPWR _21016_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23840__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25064__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17007__B2 _17022_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22967_ _15463_/X _22966_/X _22251_/X _15830_/A _22576_/A VGND VGND VPWR VPWR _22968_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20011__B1 _23666_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12720_ _12716_/A _12714_/B _12720_/C VGND VGND VPWR VPWR _12720_/X sky130_fd_sc_hd__and3_4
X_24706_ _24706_/CLK _15011_/Y HRESETn VGND VGND VPWR VPWR _24706_/Q sky130_fd_sc_hd__dfrtp_4
X_21918_ _20980_/A _21916_/X _21917_/X VGND VGND VPWR VPWR _21918_/X sky130_fd_sc_hd__and3_4
XFILLER_55_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22898_ _21030_/X _22897_/X _22646_/X _24422_/Q _22647_/X VGND VGND VPWR VPWR _22898_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12651_ _12593_/Y _12737_/A _12651_/C _12651_/D VGND VGND VPWR VPWR _12651_/X sky130_fd_sc_hd__or4_4
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24637_ _23762_/CLK _15265_/X HRESETn VGND VGND VPWR VPWR _24637_/Q sky130_fd_sc_hd__dfrtp_4
X_21849_ _21042_/A _21848_/X _22197_/A _25195_/Q _22198_/A VGND VGND VPWR VPWR _21849_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_70_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _11533_/X _15920_/A _15788_/A _25200_/Q _11537_/X VGND VGND VPWR VPWR _25200_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_30_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ _12582_/A VGND VGND VPWR VPWR _12582_/Y sky130_fd_sc_hd__inv_2
X_15370_ _15368_/X _15319_/Y _15369_/X _24598_/Q _15325_/A VGND VGND VPWR VPWR _24598_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21511__B1 _21242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24568_ _24545_/CLK _15485_/X HRESETn VGND VGND VPWR VPWR _24568_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14321_ _14319_/X _14320_/Y _24780_/Q VGND VGND VPWR VPWR _14321_/X sky130_fd_sc_hd__a21o_4
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ _11532_/X VGND VGND VPWR VPWR _11533_/X sky130_fd_sc_hd__buf_2
XFILLER_12_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23519_ _23511_/CLK _18918_/X VGND VGND VPWR VPWR _18917_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24499_ _23949_/CLK _24499_/D HRESETn VGND VGND VPWR VPWR _24499_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ _17040_/A _17116_/A _16968_/Y _17097_/A VGND VGND VPWR VPWR _17040_/X sky130_fd_sc_hd__or4_4
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14252_ _24805_/Q VGND VGND VPWR VPWR _14252_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13203_ _13203_/A _13201_/X _13202_/X VGND VGND VPWR VPWR _13207_/B sky130_fd_sc_hd__and3_4
XANTENNA__12555__B2 _24518_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14183_ _14175_/X _14182_/X _25153_/Q _14180_/X VGND VGND VPWR VPWR _14183_/X sky130_fd_sc_hd__o22a_4
XFILLER_136_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23999__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13134_ _13011_/X _13126_/X _13133_/X VGND VGND VPWR VPWR _13134_/X sky130_fd_sc_hd__and3_4
XFILLER_48_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23928__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18991_ _18990_/Y VGND VGND VPWR VPWR _18991_/X sky130_fd_sc_hd__buf_2
XANTENNA__24806__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13065_ _13075_/A VGND VGND VPWR VPWR _13065_/X sky130_fd_sc_hd__buf_2
X_17942_ _14577_/X _23439_/Q VGND VGND VPWR VPWR _17942_/X sky130_fd_sc_hd__or2_4
XANTENNA__24869__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21578__B1 _20800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12016_ _12016_/A _12016_/B VGND VGND VPWR VPWR _12016_/X sky130_fd_sc_hd__and2_4
XFILLER_78_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17873_ _17969_/A _17873_/B _17872_/X VGND VGND VPWR VPWR _17873_/X sky130_fd_sc_hd__or3_4
XFILLER_120_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16824_ _16824_/A VGND VGND VPWR VPWR _16826_/C sky130_fd_sc_hd__inv_2
X_19612_ _23273_/Q VGND VGND VPWR VPWR _21336_/B sky130_fd_sc_hd__inv_2
XFILLER_78_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22790__A2 _22788_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19543_ _19543_/A VGND VGND VPWR VPWR _21462_/B sky130_fd_sc_hd__inv_2
X_16755_ _15844_/Y _24084_/Q _15844_/Y _24084_/Q VGND VGND VPWR VPWR _16756_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13967_ _13967_/A VGND VGND VPWR VPWR _13967_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15706_ _11630_/A VGND VGND VPWR VPWR _15706_/X sky130_fd_sc_hd__buf_2
XANTENNA__24787__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12918_ _12920_/B VGND VGND VPWR VPWR _12919_/B sky130_fd_sc_hd__inv_2
X_19474_ _19472_/Y _19468_/X _19424_/X _19473_/X VGND VGND VPWR VPWR _19474_/X sky130_fd_sc_hd__a2bb2o_4
X_16686_ _24366_/Q _16685_/Y _15933_/Y _16693_/A VGND VGND VPWR VPWR _16686_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13898_ _13898_/A _13898_/B _13878_/D _13842_/X VGND VGND VPWR VPWR _13899_/B sky130_fd_sc_hd__or4_4
X_18425_ _18425_/A _18535_/A VGND VGND VPWR VPWR _18426_/D sky130_fd_sc_hd__or2_4
XANTENNA__24716__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15637_ _13612_/A _24616_/Q _14013_/A VGND VGND VPWR VPWR _15637_/X sky130_fd_sc_hd__or3_4
X_12849_ _22913_/A VGND VGND VPWR VPWR _12849_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_2_0_HCLK_A clkbuf_5_2_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15350__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18356_ _16473_/Y _18355_/X _16473_/Y _18355_/X VGND VGND VPWR VPWR _18356_/X sky130_fd_sc_hd__a2bb2o_4
X_15568_ _11527_/Y VGND VGND VPWR VPWR _20806_/A sky130_fd_sc_hd__buf_2
XANTENNA__16509__B1 _16261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22845__A3 _22459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17307_ _24001_/Q VGND VGND VPWR VPWR _17349_/A sky130_fd_sc_hd__inv_2
X_14519_ _21752_/A VGND VGND VPWR VPWR _14519_/Y sky130_fd_sc_hd__inv_2
X_18287_ _18284_/A _18277_/B _18286_/X VGND VGND VPWR VPWR _18287_/X sky130_fd_sc_hd__and3_4
X_15499_ _11585_/A VGND VGND VPWR VPWR _15499_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17238_ _17237_/Y _25221_/Q _17237_/Y _25221_/Q VGND VGND VPWR VPWR _17238_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15193__C1 _15147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17169_ _17086_/X _17160_/B _17168_/X VGND VGND VPWR VPWR _24027_/D sky130_fd_sc_hd__and3_4
XFILLER_127_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16288__A2 _16276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20180_ _23779_/Q _20234_/B VGND VGND VPWR VPWR _20189_/A sky130_fd_sc_hd__and2_4
XANTENNA__23669__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15496__B1 _24561_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23870_ _23872_/CLK _23870_/D HRESETn VGND VGND VPWR VPWR _18199_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20792__A1 _20759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20792__B2 _12062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22821_ _21572_/B _22820_/X _22640_/X _11547_/A _22641_/X VGND VGND VPWR VPWR _22821_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_42_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13673__A1_N _13446_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22752_ _16497_/Y _20807_/X VGND VGND VPWR VPWR _22752_/X sky130_fd_sc_hd__and2_4
XANTENNA__20544__B2 _20465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21741__B1 _23616_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24457__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21703_ _21694_/X _21703_/B VGND VGND VPWR VPWR _21703_/X sky130_fd_sc_hd__and2_4
X_22683_ _20643_/Y _22279_/X _20508_/A _22322_/A VGND VGND VPWR VPWR _22683_/X sky130_fd_sc_hd__o22a_4
X_21634_ _21630_/X _21633_/X _17639_/A VGND VGND VPWR VPWR _21634_/X sky130_fd_sc_hd__o21a_4
X_24422_ _24425_/CLK _24422_/D HRESETn VGND VGND VPWR VPWR _24422_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21565_ _21565_/A VGND VGND VPWR VPWR _21569_/A sky130_fd_sc_hd__buf_2
X_24353_ _24333_/CLK _16053_/X HRESETn VGND VGND VPWR VPWR _24353_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20516_ _20511_/X _20514_/X _24605_/Q _20515_/X VGND VGND VPWR VPWR _23716_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_122_0_HCLK clkbuf_7_61_0_HCLK/X VGND VGND VPWR VPWR _24333_/CLK sky130_fd_sc_hd__clkbuf_1
X_23304_ _23303_/CLK _23304_/D VGND VGND VPWR VPWR _23304_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15723__A1 _15712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24284_ _24662_/CLK _16244_/X HRESETn VGND VGND VPWR VPWR _24284_/Q sky130_fd_sc_hd__dfrtp_4
X_21496_ _13337_/A _21496_/B _21495_/X VGND VGND VPWR VPWR _21496_/X sky130_fd_sc_hd__and3_4
XFILLER_20_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_185_0_HCLK clkbuf_7_92_0_HCLK/X VGND VGND VPWR VPWR _24573_/CLK sky130_fd_sc_hd__clkbuf_1
X_23235_ _23292_/CLK _19722_/X VGND VGND VPWR VPWR _23235_/Q sky130_fd_sc_hd__dfxtp_4
X_20447_ _13506_/A VGND VGND VPWR VPWR _20447_/Y sky130_fd_sc_hd__inv_2
X_23166_ _23332_/CLK _19907_/X VGND VGND VPWR VPWR _19903_/A sky130_fd_sc_hd__dfxtp_4
X_20378_ _17179_/B _20377_/Y _20373_/X VGND VGND VPWR VPWR _20378_/X sky130_fd_sc_hd__and3_4
X_22117_ _24367_/Q _21543_/A VGND VGND VPWR VPWR _22117_/X sky130_fd_sc_hd__or2_4
XFILLER_122_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12124__A _24546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23097_ _23343_/CLK _20087_/X VGND VGND VPWR VPWR _23097_/Q sky130_fd_sc_hd__dfxtp_4
X_22048_ _22041_/Y _22046_/X _22047_/X _24932_/Q _21400_/A VGND VGND VPWR VPWR _22048_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_121_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22221__A1 _22216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11963__A _22564_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14870_ _14870_/A _15087_/A _15092_/A _14716_/Y VGND VGND VPWR VPWR _15058_/A sky130_fd_sc_hd__or4_4
XFILLER_29_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13821_ _13820_/X VGND VGND VPWR VPWR _13822_/B sky130_fd_sc_hd__inv_2
XFILLER_47_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23999_ _23992_/CLK _23999_/D HRESETn VGND VGND VPWR VPWR _17246_/A sky130_fd_sc_hd__dfrtp_4
X_16540_ _16539_/Y _16535_/X _16373_/X _16535_/X VGND VGND VPWR VPWR _24164_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24880__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13752_ _13718_/B VGND VGND VPWR VPWR _13761_/B sky130_fd_sc_hd__buf_2
XFILLER_71_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24198__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12703_ _25058_/Q _12703_/B VGND VGND VPWR VPWR _12703_/X sky130_fd_sc_hd__or2_4
X_16471_ _16471_/A VGND VGND VPWR VPWR _16471_/Y sky130_fd_sc_hd__inv_2
X_13683_ _13681_/X _13682_/Y _20201_/B VGND VGND VPWR VPWR _13683_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16266__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18210_ _18312_/A _18210_/B _18316_/A _18318_/A VGND VGND VPWR VPWR _18210_/X sky130_fd_sc_hd__or4_4
XANTENNA__24127__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15422_ _15422_/A _16475_/B VGND VGND VPWR VPWR _15422_/X sky130_fd_sc_hd__or2_4
XFILLER_31_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12634_ _12933_/C VGND VGND VPWR VPWR _12915_/C sky130_fd_sc_hd__buf_2
X_19190_ _19189_/X VGND VGND VPWR VPWR _19196_/A sky130_fd_sc_hd__inv_2
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18141_ _23866_/Q VGND VGND VPWR VPWR _18268_/A sky130_fd_sc_hd__inv_2
XFILLER_15_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15353_ _15353_/A VGND VGND VPWR VPWR _15353_/X sky130_fd_sc_hd__buf_2
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12565_ _25056_/Q VGND VGND VPWR VPWR _12565_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_81_0_HCLK clkbuf_6_40_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_81_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14304_ _16216_/A VGND VGND VPWR VPWR _14304_/X sky130_fd_sc_hd__buf_2
XFILLER_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11516_ _16231_/A _11516_/B VGND VGND VPWR VPWR _15916_/A sky130_fd_sc_hd__or2_4
X_18072_ _23896_/Q VGND VGND VPWR VPWR _18072_/X sky130_fd_sc_hd__buf_2
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15284_ _15284_/A VGND VGND VPWR VPWR _15284_/Y sky130_fd_sc_hd__inv_2
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12496_ _12495_/X VGND VGND VPWR VPWR _12497_/B sky130_fd_sc_hd__inv_2
XFILLER_8_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17023_ _24053_/Q VGND VGND VPWR VPWR _17023_/Y sky130_fd_sc_hd__inv_2
X_14235_ HWDATA[5] VGND VGND VPWR VPWR _16376_/A sky130_fd_sc_hd__buf_2
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14166_ _14160_/A _14170_/B _14145_/X VGND VGND VPWR VPWR _14166_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__15478__B1 _24571_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13117_ _13057_/X _13115_/X _25002_/Q _13116_/X VGND VGND VPWR VPWR _25002_/D sky130_fd_sc_hd__o22a_4
X_14097_ _14096_/Y _14091_/X _13645_/X _14079_/A VGND VGND VPWR VPWR _24855_/D sky130_fd_sc_hd__a2bb2o_4
X_18974_ _13123_/B VGND VGND VPWR VPWR _18974_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22450__B _12063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13048_ _18085_/A _23606_/Q VGND VGND VPWR VPWR _13048_/X sky130_fd_sc_hd__or2_4
X_17925_ _17782_/A _18800_/A VGND VGND VPWR VPWR _17926_/C sky130_fd_sc_hd__or2_4
XFILLER_100_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17856_ _17821_/A _23586_/Q VGND VGND VPWR VPWR _17857_/C sky130_fd_sc_hd__or2_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16978__B1 _16157_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16807_ _24423_/Q _16853_/A _15899_/Y _16835_/A VGND VGND VPWR VPWR _16809_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17787_ _17924_/A _18768_/A VGND VGND VPWR VPWR _17789_/B sky130_fd_sc_hd__or2_4
X_14999_ _15014_/A _14997_/X _14998_/X VGND VGND VPWR VPWR _24709_/D sky130_fd_sc_hd__and3_4
XFILLER_94_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19916__B1 _19828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16738_ _24382_/Q _17502_/B _15950_/Y _23962_/Q VGND VGND VPWR VPWR _16739_/D sky130_fd_sc_hd__a2bb2o_4
X_19526_ _19525_/Y _19523_/X _19462_/X _19523_/X VGND VGND VPWR VPWR _23304_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22178__A _22178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24550__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19457_ _19457_/A VGND VGND VPWR VPWR _19457_/Y sky130_fd_sc_hd__inv_2
X_16669_ _16652_/X _16653_/X _15704_/X _24097_/Q _16647_/X VGND VGND VPWR VPWR _24097_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_34_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15402__B1 _15286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18408_ _18378_/X _18408_/B VGND VGND VPWR VPWR _18448_/A sky130_fd_sc_hd__or2_4
XFILLER_34_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19388_ _19385_/Y _19386_/X _19387_/X _19386_/X VGND VGND VPWR VPWR _19388_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18339_ _16445_/Y _18338_/X _16445_/Y _18338_/X VGND VGND VPWR VPWR _18347_/A sky130_fd_sc_hd__a2bb2o_4
X_21350_ _21350_/A _21350_/B _21349_/X VGND VGND VPWR VPWR _21350_/X sky130_fd_sc_hd__and3_4
X_20301_ _20301_/A _20298_/A VGND VGND VPWR VPWR _20301_/Y sky130_fd_sc_hd__nand2_4
X_21281_ _21019_/A VGND VGND VPWR VPWR _21562_/A sky130_fd_sc_hd__buf_2
XFILLER_128_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13192__A1 _11711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23020_ _16389_/A _23020_/B VGND VGND VPWR VPWR _23023_/B sky130_fd_sc_hd__or2_4
X_20232_ _20232_/A _15250_/A _20232_/C VGND VGND VPWR VPWR _20232_/X sky130_fd_sc_hd__and3_4
XANTENNA__20057__A3 _13665_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22641__A _21292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15469__B1 _24575_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20163_ _20192_/A _23779_/Q _20163_/C VGND VGND VPWR VPWR _20163_/X sky130_fd_sc_hd__or3_4
XANTENNA__16130__A1 _15411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17735__A _17721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16681__A2 _13480_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21257__A _21257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20094_ _20093_/Y _20089_/X _19755_/X _20076_/Y VGND VGND VPWR VPWR _20094_/X sky130_fd_sc_hd__a2bb2o_4
X_24971_ _25186_/CLK _13483_/X HRESETn VGND VGND VPWR VPWR _13403_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12879__A _22712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23922_ _25159_/CLK _23922_/D HRESETn VGND VGND VPWR VPWR _23922_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20765__B2 _21357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16997__A2_N _24039_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24638__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23853_ _23845_/CLK _18315_/X HRESETn VGND VGND VPWR VPWR _23853_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19294__A2_N _19289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18566__A _18562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22804_ _24150_/Q _22505_/X _22576_/X _22803_/X VGND VGND VPWR VPWR _22805_/C sky130_fd_sc_hd__a211o_4
X_20996_ _21007_/A _20993_/X _20996_/C VGND VGND VPWR VPWR _20996_/X sky130_fd_sc_hd__and3_4
XFILLER_77_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23784_ _23789_/CLK _23784_/D HRESETn VGND VGND VPWR VPWR _11881_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_53_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24291__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22735_ _25092_/Q _22956_/B VGND VGND VPWR VPWR _22738_/B sky130_fd_sc_hd__or2_4
XANTENNA__24220__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22666_ _12854_/Y _20838_/X _17497_/D _22191_/X VGND VGND VPWR VPWR _22666_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22816__A _22681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21720__A _14937_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24405_ _24405_/CLK _24405_/D HRESETn VGND VGND VPWR VPWR _24405_/Q sky130_fd_sc_hd__dfrtp_4
X_21617_ _21617_/A _19606_/Y VGND VGND VPWR VPWR _21617_/X sky130_fd_sc_hd__or2_4
XFILLER_138_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19397__A _19396_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17146__B1 _17057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16814__A _17067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22597_ _22597_/A _22596_/X VGND VGND VPWR VPWR _22597_/X sky130_fd_sc_hd__and2_4
XANTENNA__22535__B _22509_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12350_ _12348_/A _12349_/A _12534_/A _12349_/Y VGND VGND VPWR VPWR _12350_/X sky130_fd_sc_hd__o22a_4
X_24336_ _24222_/CLK _24336_/D HRESETn VGND VGND VPWR VPWR _24336_/Q sky130_fd_sc_hd__dfrtp_4
X_21548_ _21540_/X _21545_/X _21546_/X _21547_/X VGND VGND VPWR VPWR _21548_/X sky130_fd_sc_hd__o22a_4
XFILLER_127_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17629__B _17629_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12281_ _12103_/Y _12281_/B VGND VGND VPWR VPWR _12281_/Y sky130_fd_sc_hd__nand2_4
X_21479_ _21346_/A _21477_/X _21478_/X VGND VGND VPWR VPWR _21479_/X sky130_fd_sc_hd__and3_4
X_24267_ _24140_/CLK _16275_/X HRESETn VGND VGND VPWR VPWR _24267_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20055__B _14197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14020_ _14020_/A _16038_/D VGND VGND VPWR VPWR _20852_/A sky130_fd_sc_hd__or2_4
X_23218_ _23112_/CLK _19770_/X VGND VGND VPWR VPWR _19769_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24198_ _24197_/CLK _16456_/X HRESETn VGND VGND VPWR VPWR _24198_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19247__A2_N _19244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23149_ _23596_/CLK _23149_/D VGND VGND VPWR VPWR _23149_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22135__A2_N _22637_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15971_ _15970_/Y _15966_/X _11594_/X _15966_/X VGND VGND VPWR VPWR _15971_/X sky130_fd_sc_hd__a2bb2o_4
X_17710_ _17674_/A VGND VGND VPWR VPWR _17889_/A sky130_fd_sc_hd__buf_2
XFILLER_96_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14922_ _24659_/Q VGND VGND VPWR VPWR _15208_/A sky130_fd_sc_hd__inv_2
X_18690_ _19303_/A _18690_/B _11734_/Y _11746_/Y VGND VGND VPWR VPWR _18690_/X sky130_fd_sc_hd__or4_4
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17641_ _17648_/B _17640_/Y _17639_/X _17648_/B VGND VGND VPWR VPWR _23940_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24379__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14853_ _15042_/A _24139_/Q _15042_/A _24139_/Q VGND VGND VPWR VPWR _14855_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15632__B1 _24505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24308__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13804_ _24903_/Q VGND VGND VPWR VPWR _13845_/A sky130_fd_sc_hd__buf_2
X_17572_ _22473_/A _17572_/B VGND VGND VPWR VPWR _17572_/X sky130_fd_sc_hd__or2_4
X_14784_ _14784_/A _14784_/B _14784_/C _14784_/D VGND VGND VPWR VPWR _14784_/X sky130_fd_sc_hd__or4_4
XFILLER_90_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11996_ _11994_/Y _11990_/X _11612_/X _11995_/X VGND VGND VPWR VPWR _11996_/X sky130_fd_sc_hd__a2bb2o_4
X_19311_ _18743_/X VGND VGND VPWR VPWR _19311_/X sky130_fd_sc_hd__buf_2
X_16523_ _16499_/A VGND VGND VPWR VPWR _16523_/X sky130_fd_sc_hd__buf_2
X_13735_ _13735_/A _13734_/Y VGND VGND VPWR VPWR _13735_/X sky130_fd_sc_hd__or2_4
XFILLER_91_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19242_ _21927_/B _19239_/X _11839_/X _19239_/X VGND VGND VPWR VPWR _19242_/X sky130_fd_sc_hd__a2bb2o_4
X_16454_ _24198_/Q VGND VGND VPWR VPWR _16454_/Y sky130_fd_sc_hd__inv_2
X_13666_ _13415_/Y _13661_/X _13665_/X _13661_/X VGND VGND VPWR VPWR _24931_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14738__A2 _14737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15405_ _24584_/Q VGND VGND VPWR VPWR _15405_/Y sky130_fd_sc_hd__inv_2
X_12617_ _24522_/Q VGND VGND VPWR VPWR _12617_/Y sky130_fd_sc_hd__inv_2
X_19173_ _19172_/Y _19169_/X _19149_/X _19169_/X VGND VGND VPWR VPWR _19173_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16385_ _24223_/Q VGND VGND VPWR VPWR _16385_/Y sky130_fd_sc_hd__inv_2
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13597_ _13559_/B _13596_/Y _13594_/X _13587_/X _11670_/A VGND VGND VPWR VPWR _13597_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18124_ _18124_/A VGND VGND VPWR VPWR _18124_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22445__B _22445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15336_ _22884_/A _15333_/X _11540_/X _15333_/X VGND VGND VPWR VPWR _24611_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18642__C _14482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12548_ _25043_/Q _12546_/Y _12547_/Y _24529_/Q VGND VGND VPWR VPWR _12552_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23943__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25167__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15699__B1 _15513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18055_ _18054_/X VGND VGND VPWR VPWR _18055_/Y sky130_fd_sc_hd__inv_2
X_15267_ _14100_/X _14074_/A _15240_/A _13745_/B _15262_/X VGND VGND VPWR VPWR _24635_/D
+ sky130_fd_sc_hd__a32o_4
X_12479_ _12412_/A _12478_/X VGND VGND VPWR VPWR _12479_/Y sky130_fd_sc_hd__nand2_4
X_17006_ _24055_/Q VGND VGND VPWR VPWR _17022_/B sky130_fd_sc_hd__inv_2
X_14218_ _14218_/A VGND VGND VPWR VPWR _14218_/X sky130_fd_sc_hd__buf_2
X_15198_ _15112_/A _15197_/X VGND VGND VPWR VPWR _15219_/A sky130_fd_sc_hd__or2_4
Xclkbuf_8_25_0_HCLK clkbuf_7_12_0_HCLK/X VGND VGND VPWR VPWR _25186_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_98_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22984__A2 _22859_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14149_ _20889_/A _12053_/A VGND VGND VPWR VPWR _14149_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_88_0_HCLK clkbuf_7_44_0_HCLK/X VGND VGND VPWR VPWR _24823_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12789__A1_N _22258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18957_ _17903_/B VGND VGND VPWR VPWR _18957_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13477__A2 _13480_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12699__A _12638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15871__B1 _11581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17908_ _17708_/X _17907_/X _23928_/Q _17767_/X VGND VGND VPWR VPWR _23928_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19062__B1 _19038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18888_ _23530_/Q VGND VGND VPWR VPWR _18888_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24731__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17839_ _17903_/A _17839_/B VGND VGND VPWR VPWR _17839_/X sky130_fd_sc_hd__or2_4
XFILLER_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15623__B1 _15511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24049__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20850_ _20850_/A VGND VGND VPWR VPWR _20850_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19509_ _19862_/A _19883_/B _19509_/C VGND VGND VPWR VPWR _19509_/X sky130_fd_sc_hd__or3_4
X_20781_ _20800_/A VGND VGND VPWR VPWR _20782_/A sky130_fd_sc_hd__buf_2
XFILLER_63_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22520_ _21978_/X _22519_/X VGND VGND VPWR VPWR _22520_/X sky130_fd_sc_hd__and2_4
XFILLER_23_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21540__A _22637_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13042__B _23134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22451_ _13609_/X _22449_/X _20902_/X _22450_/Y VGND VGND VPWR VPWR _22451_/X sky130_fd_sc_hd__o22a_4
XFILLER_10_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21402_ _21047_/A VGND VGND VPWR VPWR _21402_/X sky130_fd_sc_hd__buf_2
X_22382_ _24373_/Q _22238_/X VGND VGND VPWR VPWR _22382_/X sky130_fd_sc_hd__or2_4
XANTENNA__23684__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25170_ _23288_/CLK _25170_/D HRESETn VGND VGND VPWR VPWR _11855_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17449__B _17460_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12881__B _12947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20156__A _14206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21333_ _21333_/A _19679_/Y VGND VGND VPWR VPWR _21334_/C sky130_fd_sc_hd__or2_4
X_24121_ _24094_/CLK _24121_/D HRESETn VGND VGND VPWR VPWR _14777_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21880__C1 _21879_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21264_ _22501_/A _21263_/X _21036_/X _24547_/Q _11530_/X VGND VGND VPWR VPWR _21265_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_85_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24052_ _24049_/CLK _24052_/D HRESETn VGND VGND VPWR VPWR _17080_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_137_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20215_ _20204_/X _23773_/Q VGND VGND VPWR VPWR _20227_/A sky130_fd_sc_hd__and2_4
X_23003_ _22335_/A _23002_/X _22835_/X _25221_/Q _22576_/A VGND VGND VPWR VPWR _23003_/X
+ sky130_fd_sc_hd__a32o_4
X_21195_ _21008_/A VGND VGND VPWR VPWR _21238_/A sky130_fd_sc_hd__buf_2
XANTENNA__18596__A1_N _24243_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20146_ _20145_/Y _20141_/X _15522_/X _20141_/X VGND VGND VPWR VPWR _23072_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24819__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22727__A2 _21544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19680__A _19680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20077_ _20076_/Y VGND VGND VPWR VPWR _20077_/X sky130_fd_sc_hd__buf_2
X_24954_ _24824_/CLK _24954_/D HRESETn VGND VGND VPWR VPWR _24954_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12402__A _12451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24472__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23905_ _24937_/CLK _23905_/D HRESETn VGND VGND VPWR VPWR _23040_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_72_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24885_ _24884_/CLK _24885_/D HRESETn VGND VGND VPWR VPWR _13926_/C sky130_fd_sc_hd__dfrtp_4
XANTENNA__15614__B1 _24517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24401__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11850_ _11850_/A VGND VGND VPWR VPWR _19614_/A sky130_fd_sc_hd__buf_2
X_23836_ _23828_/CLK _18480_/X HRESETn VGND VGND VPWR VPWR _18388_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_61_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14233__A1_N _14230_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11781_ _11694_/X VGND VGND VPWR VPWR _13551_/B sky130_fd_sc_hd__inv_2
X_23767_ _23767_/CLK _20260_/X HRESETn VGND VGND VPWR VPWR _23767_/Q sky130_fd_sc_hd__dfrtp_4
X_20979_ _20979_/A _19300_/Y VGND VGND VPWR VPWR _20980_/C sky130_fd_sc_hd__or2_4
XFILLER_82_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13520_ _20740_/A _13518_/X _13519_/Y VGND VGND VPWR VPWR _13520_/X sky130_fd_sc_hd__o21a_4
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15917__A1 _11535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22718_ _22718_/A _22699_/X _22661_/C _22718_/D VGND VGND VPWR VPWR HRDATA[21] sky130_fd_sc_hd__or4_4
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23698_ _24349_/CLK _23698_/D HRESETn VGND VGND VPWR VPWR _23698_/Q sky130_fd_sc_hd__dfrtp_4
X_13451_ _13449_/A VGND VGND VPWR VPWR _14394_/A sky130_fd_sc_hd__inv_2
X_22649_ _22637_/X _22643_/Y _22601_/X _22648_/X VGND VGND VPWR VPWR _22649_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22265__B _22265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12402_ _12451_/A _12448_/A VGND VGND VPWR VPWR _12402_/X sky130_fd_sc_hd__or2_4
X_16170_ _16165_/A VGND VGND VPWR VPWR _16170_/X sky130_fd_sc_hd__buf_2
XANTENNA__22663__A1 _12617_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13382_ _13381_/Y _13377_/X _13330_/X _13377_/X VGND VGND VPWR VPWR _24977_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22663__B2 _22029_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15121_ _14885_/Y _15118_/X VGND VGND VPWR VPWR _15121_/X sky130_fd_sc_hd__or2_4
X_12333_ _25094_/Q _24491_/Q _12448_/A _12332_/Y VGND VGND VPWR VPWR _12337_/C sky130_fd_sc_hd__o22a_4
X_24319_ _24319_/CLK _24319_/D HRESETn VGND VGND VPWR VPWR _24319_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15052_ _24695_/Q _15051_/Y VGND VGND VPWR VPWR _15052_/X sky130_fd_sc_hd__or2_4
X_12264_ _12091_/Y _12167_/Y VGND VGND VPWR VPWR _12298_/A sky130_fd_sc_hd__or2_4
XANTENNA__22281__A _20900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_241_0_HCLK clkbuf_8_241_0_HCLK/A VGND VGND VPWR VPWR _24145_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_123_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14003_ _14002_/X VGND VGND VPWR VPWR _14003_/Y sky130_fd_sc_hd__inv_2
X_12195_ _12538_/B VGND VGND VPWR VPWR _12195_/X sky130_fd_sc_hd__buf_2
X_19860_ _21002_/B _19854_/X _19859_/X _19841_/X VGND VGND VPWR VPWR _19860_/X sky130_fd_sc_hd__a2bb2o_4
X_18811_ _13061_/B VGND VGND VPWR VPWR _18811_/Y sky130_fd_sc_hd__inv_2
X_19791_ _21522_/B _19786_/X _19455_/X _19786_/X VGND VGND VPWR VPWR _23210_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22179__B1 _12329_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15954_ _15952_/Y _15948_/X _15772_/X _15953_/X VGND VGND VPWR VPWR _15954_/X sky130_fd_sc_hd__a2bb2o_4
X_18742_ _18742_/A VGND VGND VPWR VPWR _18742_/Y sky130_fd_sc_hd__inv_2
X_14905_ _14896_/X _14905_/B _14905_/C _14904_/X VGND VGND VPWR VPWR _14932_/B sky130_fd_sc_hd__or4_4
X_18673_ _18682_/A VGND VGND VPWR VPWR _18673_/X sky130_fd_sc_hd__buf_2
X_15885_ _15885_/A VGND VGND VPWR VPWR _15885_/X sky130_fd_sc_hd__buf_2
XFILLER_64_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15605__B1 _15350_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24142__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14836_ _14836_/A VGND VGND VPWR VPWR _14836_/Y sky130_fd_sc_hd__inv_2
X_17624_ _17460_/B VGND VGND VPWR VPWR _17625_/A sky130_fd_sc_hd__buf_2
XFILLER_5_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17555_ _17547_/X _17553_/X _17554_/X VGND VGND VPWR VPWR _17555_/X sky130_fd_sc_hd__and3_4
XANTENNA__15620__A3 _15507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14767_ _15004_/A _24116_/Q _14765_/Y _24116_/Q VGND VGND VPWR VPWR _14773_/B sky130_fd_sc_hd__a2bb2o_4
X_11979_ _11977_/Y _11978_/X _11636_/X _11978_/X VGND VGND VPWR VPWR _25150_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14239__A _24812_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16506_ _16499_/A VGND VGND VPWR VPWR _16506_/X sky130_fd_sc_hd__buf_2
X_13718_ _13753_/C _13718_/B _13766_/D VGND VGND VPWR VPWR _13718_/X sky130_fd_sc_hd__or3_4
X_17486_ _17486_/A _21839_/A VGND VGND VPWR VPWR _17486_/X sky130_fd_sc_hd__or2_4
X_14698_ _14697_/Y _24124_/Q _14697_/Y _24124_/Q VGND VGND VPWR VPWR _14698_/X sky130_fd_sc_hd__a2bb2o_4
X_16437_ _16436_/Y _16434_/X _16087_/X _16434_/X VGND VGND VPWR VPWR _16437_/X sky130_fd_sc_hd__a2bb2o_4
X_19225_ _19225_/A VGND VGND VPWR VPWR _19225_/Y sky130_fd_sc_hd__inv_2
X_13649_ _13649_/A VGND VGND VPWR VPWR _13649_/X sky130_fd_sc_hd__buf_2
XFILLER_20_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22027__A2_N _21544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19156_ _19155_/Y _19153_/X _19109_/X _19153_/X VGND VGND VPWR VPWR _23435_/D sky130_fd_sc_hd__a2bb2o_4
X_16368_ _24229_/Q VGND VGND VPWR VPWR _16368_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18107_ _18095_/X _18093_/Y _18106_/X _21644_/A _18096_/Y VGND VGND VPWR VPWR _23887_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_121_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_51_0_HCLK clkbuf_6_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_51_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_15319_ _15531_/B VGND VGND VPWR VPWR _15319_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11598__A _16100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19087_ _19086_/Y _19084_/X _18953_/X _19084_/X VGND VGND VPWR VPWR _23459_/D sky130_fd_sc_hd__a2bb2o_4
X_16299_ _21882_/A VGND VGND VPWR VPWR _16300_/A sky130_fd_sc_hd__buf_2
X_18038_ _18038_/A _17460_/B VGND VGND VPWR VPWR _18038_/X sky130_fd_sc_hd__or2_4
XANTENNA__15687__A3 _16087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22191__A _11516_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24983__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20000_ _20000_/A VGND VGND VPWR VPWR _20000_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16097__B1 _16096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24912__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19989_ _11755_/A _18075_/X _11734_/Y _18064_/X VGND VGND VPWR VPWR _19989_/X sky130_fd_sc_hd__or4_4
XFILLER_45_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21951_ _21394_/A _21951_/B _21950_/X VGND VGND VPWR VPWR _21951_/X sky130_fd_sc_hd__and3_4
X_20902_ _11720_/X VGND VGND VPWR VPWR _20902_/X sky130_fd_sc_hd__buf_2
X_24670_ _24671_/CLK _24670_/D HRESETn VGND VGND VPWR VPWR _24670_/Q sky130_fd_sc_hd__dfrtp_4
X_21882_ _21882_/A VGND VGND VPWR VPWR _21882_/X sky130_fd_sc_hd__buf_2
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _24769_/CLK _20716_/X HRESETn VGND VGND VPWR VPWR _13863_/A sky130_fd_sc_hd__dfrtp_4
X_20833_ _22858_/A VGND VGND VPWR VPWR _20833_/X sky130_fd_sc_hd__buf_2
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16967__A1_N _16193_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14149__A _20889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23865__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23552_ _23537_/CLK _18826_/X VGND VGND VPWR VPWR _13258_/B sky130_fd_sc_hd__dfxtp_4
X_20764_ _22014_/B _20762_/X _24321_/Q _21591_/B VGND VGND VPWR VPWR _20764_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22366__A _22198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25089__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22503_ _24271_/Q _22350_/X _22351_/X VGND VGND VPWR VPWR _22503_/X sky130_fd_sc_hd__o21a_4
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20695_ _12026_/X _20695_/B VGND VGND VPWR VPWR _20695_/X sky130_fd_sc_hd__and2_4
XFILLER_56_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23483_ _23482_/CLK _19021_/X VGND VGND VPWR VPWR _23483_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25018__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22434_ _22434_/A _20749_/X VGND VGND VPWR VPWR _22434_/X sky130_fd_sc_hd__or2_4
XFILLER_136_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25153_ _24824_/CLK _11972_/X HRESETn VGND VGND VPWR VPWR _25153_/Q sky130_fd_sc_hd__dfrtp_4
X_22365_ _22365_/A _21979_/X VGND VGND VPWR VPWR _22365_/X sky130_fd_sc_hd__or2_4
XFILLER_87_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24104_ _24104_/CLK _16660_/X HRESETn VGND VGND VPWR VPWR _16658_/A sky130_fd_sc_hd__dfrtp_4
X_21316_ _15284_/Y _11501_/X _14090_/A _20758_/X VGND VGND VPWR VPWR _21316_/X sky130_fd_sc_hd__a2bb2o_4
X_22296_ _21991_/X _22295_/X VGND VGND VPWR VPWR _22296_/X sky130_fd_sc_hd__and2_4
X_25084_ _25084_/CLK _25084_/D HRESETn VGND VGND VPWR VPWR _12362_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_11_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22948__A2 _21544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14886__B2 _24286_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21247_ _21218_/X _21244_/X _21246_/X VGND VGND VPWR VPWR _21247_/Y sky130_fd_sc_hd__a21oi_4
X_24035_ _24596_/CLK _24035_/D HRESETn VGND VGND VPWR VPWR _22164_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16088__B1 _16087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24653__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21178_ _21178_/A VGND VGND VPWR VPWR _22806_/B sky130_fd_sc_hd__buf_2
XFILLER_46_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11955__B _11954_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_71_0_HCLK clkbuf_8_71_0_HCLK/A VGND VGND VPWR VPWR _24811_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15835__B1 _15753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20129_ _17982_/A _20119_/X _11643_/A _23078_/Q _20116_/X VGND VGND VPWR VPWR _23078_/D
+ sky130_fd_sc_hd__a32o_4
X_12951_ _12951_/A _12951_/B VGND VGND VPWR VPWR _12952_/C sky130_fd_sc_hd__or2_4
XFILLER_46_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24937_ _24937_/CLK _24937_/D HRESETn VGND VGND VPWR VPWR _13411_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_46_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11971__A _11965_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11902_ _11902_/A _11893_/X _11902_/C _11901_/X VGND VGND VPWR VPWR _11902_/X sky130_fd_sc_hd__or4_4
XANTENNA__15443__A _14436_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15670_ _12320_/Y _15666_/X _11540_/X _15669_/X VGND VGND VPWR VPWR _24494_/D sky130_fd_sc_hd__a2bb2o_4
X_12882_ _12836_/Y _12829_/Y _12882_/C _12881_/X VGND VGND VPWR VPWR _12883_/B sky130_fd_sc_hd__or4_4
X_24868_ _24870_/CLK _14056_/X HRESETn VGND VGND VPWR VPWR _14055_/A sky130_fd_sc_hd__dfstp_4
XFILLER_22_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16260__B1 _16259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14621_ _14620_/Y VGND VGND VPWR VPWR _14621_/X sky130_fd_sc_hd__buf_2
X_11833_ _19714_/A VGND VGND VPWR VPWR _19600_/A sky130_fd_sc_hd__buf_2
XFILLER_33_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23819_ _23824_/CLK _23819_/D HRESETn VGND VGND VPWR VPWR _23819_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ _24788_/CLK _14269_/X HRESETn VGND VGND VPWR VPWR _13921_/A sky130_fd_sc_hd__dfrtp_4
X_17340_ _17340_/A _17339_/X VGND VGND VPWR VPWR _17340_/X sky130_fd_sc_hd__or2_4
XFILLER_57_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _17806_/A VGND VGND VPWR VPWR _17739_/A sky130_fd_sc_hd__buf_2
XPHY_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11763_/A VGND VGND VPWR VPWR _11765_/A sky130_fd_sc_hd__inv_2
XPHY_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _13503_/A _13503_/B VGND VGND VPWR VPWR _13503_/X sky130_fd_sc_hd__or2_4
XANTENNA__21180__A _21400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _25207_/Q _17270_/Y _11618_/Y _17430_/A VGND VGND VPWR VPWR _17277_/A sky130_fd_sc_hd__a2bb2o_4
X_14483_ _14476_/Y _14482_/X _21534_/A VGND VGND VPWR VPWR _14506_/B sky130_fd_sc_hd__and3_4
XFILLER_70_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _11649_/Y _11694_/X VGND VGND VPWR VPWR _11718_/B sky130_fd_sc_hd__or2_4
XFILLER_105_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19010_ _14548_/A _24739_/Q _14482_/X VGND VGND VPWR VPWR _19509_/C sky130_fd_sc_hd__or3_4
XPHY_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16222_ _16003_/Y _14431_/A _16222_/C _14435_/D VGND VGND VPWR VPWR _16223_/A sky130_fd_sc_hd__or4_4
XPHY_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13434_ _24932_/Q VGND VGND VPWR VPWR _13434_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21439__A2 _20751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14506__B _14506_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16153_ HWDATA[26] VGND VGND VPWR VPWR _16153_/X sky130_fd_sc_hd__buf_2
X_13365_ _11904_/Y _13363_/X _11607_/X _13363_/X VGND VGND VPWR VPWR _24985_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_6_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12307__A _24473_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15104_ _24671_/Q VGND VGND VPWR VPWR _15104_/Y sky130_fd_sc_hd__inv_2
X_12316_ _24477_/Q VGND VGND VPWR VPWR _12316_/Y sky130_fd_sc_hd__inv_2
X_16084_ _16084_/A VGND VGND VPWR VPWR _16084_/X sky130_fd_sc_hd__buf_2
X_13296_ _13232_/A _13292_/X _13296_/C VGND VGND VPWR VPWR _13304_/B sky130_fd_sc_hd__or3_4
X_15035_ _15035_/A _15034_/X VGND VGND VPWR VPWR _15035_/Y sky130_fd_sc_hd__nand2_4
X_19912_ _21787_/B _19906_/X _19821_/X _19911_/X VGND VGND VPWR VPWR _23164_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12247_ _12227_/X _12244_/B _12246_/Y VGND VGND VPWR VPWR _12247_/X sky130_fd_sc_hd__and3_4
XFILLER_64_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16079__B1 _15775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24394__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19843_ _22057_/B _19842_/X _19815_/X _19842_/X VGND VGND VPWR VPWR _23190_/D sky130_fd_sc_hd__a2bb2o_4
X_12178_ _12265_/A _12265_/B _12178_/C _12275_/A VGND VGND VPWR VPWR _12178_/X sky130_fd_sc_hd__or4_4
XFILLER_68_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11560__B1 _11558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24323__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19774_ _19774_/A VGND VGND VPWR VPWR _19774_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16986_ _16986_/A VGND VGND VPWR VPWR _17034_/A sky130_fd_sc_hd__inv_2
X_18725_ _18723_/Y _18719_/X _18679_/X _18724_/X VGND VGND VPWR VPWR _18725_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21355__A _17636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15937_ _15935_/Y _15936_/X _11545_/X _15936_/X VGND VGND VPWR VPWR _15937_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15868_ _15885_/A VGND VGND VPWR VPWR _15868_/X sky130_fd_sc_hd__buf_2
X_18656_ _23609_/Q VGND VGND VPWR VPWR _21377_/B sky130_fd_sc_hd__inv_2
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14819_ _24684_/Q _14818_/A _15087_/A _14818_/Y VGND VGND VPWR VPWR _14819_/X sky130_fd_sc_hd__o22a_4
X_17607_ _17603_/A _17607_/B _17606_/Y VGND VGND VPWR VPWR _17607_/X sky130_fd_sc_hd__and3_4
X_15799_ _16581_/A VGND VGND VPWR VPWR _15799_/X sky130_fd_sc_hd__buf_2
X_18587_ _18583_/X _18587_/B _18585_/X _18587_/D VGND VGND VPWR VPWR _18587_/X sky130_fd_sc_hd__or4_4
XFILLER_91_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17538_ _17509_/A _17538_/B _17537_/X VGND VGND VPWR VPWR _23967_/D sky130_fd_sc_hd__and3_4
XFILLER_60_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22186__A _21569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25182__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17469_ _17465_/Y _17468_/Y _17465_/A _17468_/A VGND VGND VPWR VPWR _17469_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25111__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19208_ _19206_/Y _19204_/X _19207_/X _19204_/X VGND VGND VPWR VPWR _23416_/D sky130_fd_sc_hd__a2bb2o_4
X_20480_ _13509_/B VGND VGND VPWR VPWR _20480_/Y sky130_fd_sc_hd__inv_2
X_19139_ _23440_/Q VGND VGND VPWR VPWR _19139_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14708__A1_N _15033_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22150_ _24133_/Q _22147_/X _22148_/X _22149_/X VGND VGND VPWR VPWR _22150_/X sky130_fd_sc_hd__a211o_4
XFILLER_133_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21101_ _16471_/Y _16300_/A _22858_/A VGND VGND VPWR VPWR _21101_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16719__A2_N _17558_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22081_ _14523_/A _22077_/X _22080_/X VGND VGND VPWR VPWR _22082_/C sky130_fd_sc_hd__or3_4
XFILLER_86_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21032_ _12356_/A _21408_/B VGND VGND VPWR VPWR _21032_/X sky130_fd_sc_hd__or2_4
XANTENNA__21063__B1 _21062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11775__B _11694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15817__B1 _15712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_58_0_HCLK clkbuf_7_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_58_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24064__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19008__B1 _18662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21366__A1 _21356_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22983_ _24123_/Q _22857_/B VGND VGND VPWR VPWR _22983_/X sky130_fd_sc_hd__or2_4
XFILLER_55_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24722_ _24723_/CLK _14666_/X HRESETn VGND VGND VPWR VPWR _14626_/A sky130_fd_sc_hd__dfrtp_4
X_21934_ _21158_/A _21934_/B VGND VGND VPWR VPWR _21934_/X sky130_fd_sc_hd__or2_4
XFILLER_28_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24653_ _24654_/CLK _24653_/D HRESETn VGND VGND VPWR VPWR _14964_/A sky130_fd_sc_hd__dfrtp_4
X_21865_ _21864_/X VGND VGND VPWR VPWR _21870_/A sky130_fd_sc_hd__buf_2
XANTENNA__21118__A1 _12054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ _24005_/CLK _18674_/X VGND VGND VPWR VPWR _23604_/Q sky130_fd_sc_hd__dfxtp_4
X_20816_ _12322_/A _22429_/B _20815_/X VGND VGND VPWR VPWR _20816_/X sky130_fd_sc_hd__o21a_4
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24584_ _24587_/CLK _15406_/X HRESETn VGND VGND VPWR VPWR _24584_/Q sky130_fd_sc_hd__dfrtp_4
X_21796_ _20058_/Y _21113_/B _21582_/X _21795_/Y VGND VGND VPWR VPWR _21796_/X sky130_fd_sc_hd__a211o_4
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23535_ _24998_/CLK _18871_/X VGND VGND VPWR VPWR _18870_/A sky130_fd_sc_hd__dfxtp_4
X_20747_ _15821_/X VGND VGND VPWR VPWR _20747_/X sky130_fd_sc_hd__buf_2
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14607__A scl_oen_o_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22618__A1 _24144_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23466_ _23416_/CLK _23466_/D VGND VGND VPWR VPWR _17848_/B sky130_fd_sc_hd__dfxtp_4
X_20678_ _20556_/X _20677_/X _24187_/Q _20602_/X VGND VGND VPWR VPWR _23756_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25205_ _24372_/CLK _11582_/X HRESETn VGND VGND VPWR VPWR _11579_/A sky130_fd_sc_hd__dfrtp_4
X_22417_ _22394_/X _22398_/X _22404_/Y _22416_/X VGND VGND VPWR VPWR HRDATA[13] sky130_fd_sc_hd__a211o_4
XFILLER_13_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17918__A _17918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23397_ _25194_/CLK _23397_/D VGND VGND VPWR VPWR _19263_/A sky130_fd_sc_hd__dfxtp_4
X_13150_ _11753_/A _13150_/B _13150_/C VGND VGND VPWR VPWR _13151_/C sky130_fd_sc_hd__and3_4
XANTENNA__24834__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25136_ _23796_/CLK _25136_/D HRESETn VGND VGND VPWR VPWR SCLK_S3 sky130_fd_sc_hd__dfstp_4
X_22348_ _23023_/A VGND VGND VPWR VPWR _22348_/X sky130_fd_sc_hd__buf_2
XFILLER_136_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12101_ _24569_/Q VGND VGND VPWR VPWR _12101_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11966__A _11965_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23043__A1 _22263_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13081_ _11751_/X VGND VGND VPWR VPWR _13171_/A sky130_fd_sc_hd__buf_2
X_25067_ _25067_/CLK _25067_/D HRESETn VGND VGND VPWR VPWR _25067_/Q sky130_fd_sc_hd__dfrtp_4
X_22279_ _22279_/A VGND VGND VPWR VPWR _22279_/X sky130_fd_sc_hd__buf_2
X_12032_ _25144_/Q _12031_/Y _25144_/Q _12031_/Y VGND VGND VPWR VPWR _12033_/D sky130_fd_sc_hd__a2bb2o_4
X_24018_ _23852_/CLK _17203_/X HRESETn VGND VGND VPWR VPWR _24018_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16840_ _16840_/A _16840_/B VGND VGND VPWR VPWR _16841_/D sky130_fd_sc_hd__or2_4
XANTENNA__21175__A _20777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16771_ _16771_/A VGND VGND VPWR VPWR _16771_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13983_ _13927_/A _13927_/B _13927_/A _13927_/B VGND VGND VPWR VPWR _13983_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15722_ _15717_/A _15717_/B _15722_/C VGND VGND VPWR VPWR _15722_/X sky130_fd_sc_hd__or3_4
X_18510_ _18430_/Y _18508_/A VGND VGND VPWR VPWR _18511_/C sky130_fd_sc_hd__or2_4
X_12934_ _12880_/A _12833_/X _12955_/B VGND VGND VPWR VPWR _12943_/D sky130_fd_sc_hd__or3_4
X_19490_ _19486_/Y _19489_/X _19442_/X _19489_/X VGND VGND VPWR VPWR _23318_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23787__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15653_ _21092_/B VGND VGND VPWR VPWR _15653_/X sky130_fd_sc_hd__buf_2
X_18441_ _18440_/X VGND VGND VPWR VPWR _18442_/B sky130_fd_sc_hd__inv_2
X_12865_ _12859_/X _12865_/B _12865_/C _12864_/X VGND VGND VPWR VPWR _12865_/X sky130_fd_sc_hd__or4_4
XANTENNA__23716__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15587__A2 _15582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18484__A _18484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14604_ _18873_/B VGND VGND VPWR VPWR _18759_/B sky130_fd_sc_hd__buf_2
X_11816_ _11780_/Y _11818_/A _11815_/X VGND VGND VPWR VPWR _11816_/Y sky130_fd_sc_hd__o21ai_4
X_18372_ _23822_/Q VGND VGND VPWR VPWR _18373_/A sky130_fd_sc_hd__inv_2
X_15584_ _15584_/A VGND VGND VPWR VPWR _15585_/A sky130_fd_sc_hd__buf_2
X_12796_ _22605_/A VGND VGND VPWR VPWR _12796_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17323_ _17273_/Y _17321_/Y _17323_/C _17323_/D VGND VGND VPWR VPWR _17324_/C sky130_fd_sc_hd__or4_4
XANTENNA__20868__B1 _20866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _21205_/A VGND VGND VPWR VPWR _21378_/A sky130_fd_sc_hd__buf_2
XPHY_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11746_/Y VGND VGND VPWR VPWR _11761_/A sky130_fd_sc_hd__buf_2
XPHY_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17254_ _25198_/Q _17253_/A _11606_/Y _17413_/A VGND VGND VPWR VPWR _17259_/B sky130_fd_sc_hd__o22a_4
XANTENNA__22609__A1 _23960_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466_ _14448_/X _14453_/X _14463_/Y _14465_/X VGND VGND VPWR VPWR _14466_/X sky130_fd_sc_hd__or4_4
XFILLER_105_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _11676_/A _11677_/A _11676_/Y _11677_/Y VGND VGND VPWR VPWR _11682_/C sky130_fd_sc_hd__o22a_4
XFILLER_70_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22734__A _22677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16205_ _24294_/Q VGND VGND VPWR VPWR _16205_/Y sky130_fd_sc_hd__inv_2
X_13417_ _13415_/Y _13413_/A _13655_/A _14385_/A VGND VGND VPWR VPWR _13418_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17185_ _17184_/Y VGND VGND VPWR VPWR _17185_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14397_ _14387_/A _14386_/Y VGND VGND VPWR VPWR _14397_/X sky130_fd_sc_hd__or2_4
XFILLER_128_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16136_ _16135_/X VGND VGND VPWR VPWR _16137_/A sky130_fd_sc_hd__buf_2
XANTENNA__24575__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13348_ _13348_/A VGND VGND VPWR VPWR _13348_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24504__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16067_ _16066_/Y _16064_/X _11555_/X _16064_/X VGND VGND VPWR VPWR _16067_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13279_ _13073_/A _13279_/B _13278_/X VGND VGND VPWR VPWR _13279_/X sky130_fd_sc_hd__or3_4
XANTENNA__14252__A _24805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15018_ _14867_/A VGND VGND VPWR VPWR _15018_/X sky130_fd_sc_hd__buf_2
XFILLER_116_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22793__B1 _16063_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19826_ _19824_/Y _19822_/X _19825_/X _19822_/X VGND VGND VPWR VPWR _23195_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16472__B1 _16216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19757_ _19757_/A VGND VGND VPWR VPWR _22095_/B sky130_fd_sc_hd__inv_2
XFILLER_110_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16969_ _24054_/Q VGND VGND VPWR VPWR _17070_/A sky130_fd_sc_hd__inv_2
XFILLER_84_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22545__B1 _13362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16179__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18708_ _13266_/B VGND VGND VPWR VPWR _18708_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19410__B1 _19387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19688_ _19688_/A VGND VGND VPWR VPWR _19688_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18639_ _11645_/X _18636_/X _18638_/X VGND VGND VPWR VPWR _18639_/X sky130_fd_sc_hd__o21a_4
XFILLER_25_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16775__A1 _24424_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16775__B2 _16774_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21650_ _21646_/Y _21647_/X _21648_/X _21649_/X VGND VGND VPWR VPWR _21651_/B sky130_fd_sc_hd__a211o_4
X_20601_ _20601_/A VGND VGND VPWR VPWR _20651_/A sky130_fd_sc_hd__inv_2
X_21581_ _21581_/A _12061_/B _21580_/X VGND VGND VPWR VPWR _21581_/X sky130_fd_sc_hd__and3_4
XFILLER_21_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23320_ _23336_/CLK _23320_/D VGND VGND VPWR VPWR _13284_/B sky130_fd_sc_hd__dfxtp_4
X_20532_ _13512_/C _20528_/X _20531_/Y VGND VGND VPWR VPWR _20532_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_21_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22644__A _22249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20463_ _23705_/Q _13506_/X _20462_/Y VGND VGND VPWR VPWR _20463_/Y sky130_fd_sc_hd__a21oi_4
X_23251_ _23242_/CLK _23251_/D VGND VGND VPWR VPWR _23251_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_4_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22202_ _22202_/A _22438_/A VGND VGND VPWR VPWR _22202_/X sky130_fd_sc_hd__and2_4
Xclkbuf_5_21_0_HCLK clkbuf_4_10_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20394_ _20394_/A VGND VGND VPWR VPWR _20394_/Y sky130_fd_sc_hd__inv_2
X_23182_ _23156_/CLK _23182_/D VGND VGND VPWR VPWR _23182_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24245__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22133_ _22133_/A _22527_/B VGND VGND VPWR VPWR _22133_/X sky130_fd_sc_hd__and2_4
XFILLER_121_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22064_ _22064_/A _22064_/B VGND VGND VPWR VPWR _22065_/C sky130_fd_sc_hd__or2_4
XFILLER_47_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22784__B1 _20801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21015_ _20998_/A _19527_/Y _21007_/A VGND VGND VPWR VPWR _21015_/X sky130_fd_sc_hd__o21a_4
XFILLER_88_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21707__B _21707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16463__B1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23880__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_145_0_HCLK clkbuf_7_72_0_HCLK/X VGND VGND VPWR VPWR _23993_/CLK sky130_fd_sc_hd__clkbuf_1
X_22966_ _24319_/Q _22999_/B VGND VGND VPWR VPWR _22966_/X sky130_fd_sc_hd__or2_4
XANTENNA__20011__A1 _23126_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24705_ _24671_/CLK _24705_/D HRESETn VGND VGND VPWR VPWR _24705_/Q sky130_fd_sc_hd__dfrtp_4
X_21917_ _21913_/A _21917_/B VGND VGND VPWR VPWR _21917_/X sky130_fd_sc_hd__or2_4
XFILLER_82_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16766__A1 _24414_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22897_ _24316_/Q _22897_/B VGND VGND VPWR VPWR _22897_/X sky130_fd_sc_hd__or2_4
XANTENNA__25033__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12650_ _12650_/A VGND VGND VPWR VPWR _12651_/C sky130_fd_sc_hd__inv_2
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24636_ _23762_/CLK _24636_/D HRESETn VGND VGND VPWR VPWR _13722_/A sky130_fd_sc_hd__dfrtp_4
X_21848_ _24365_/Q _21848_/B VGND VGND VPWR VPWR _21848_/X sky130_fd_sc_hd__or2_4
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ HWDATA[10] VGND VGND VPWR VPWR _15788_/A sky130_fd_sc_hd__buf_2
XANTENNA__19704__B2 _19701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ _12581_/A VGND VGND VPWR VPWR _12581_/Y sky130_fd_sc_hd__inv_2
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24567_ _24573_/CLK _15486_/X HRESETn VGND VGND VPWR VPWR _24567_/Q sky130_fd_sc_hd__dfrtp_4
X_21779_ _21519_/A _21777_/X _21779_/C VGND VGND VPWR VPWR _21779_/X sky130_fd_sc_hd__and3_4
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14320_ _23649_/Q VGND VGND VPWR VPWR _14320_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13241__A _13136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11532_ _11532_/A VGND VGND VPWR VPWR _11532_/X sky130_fd_sc_hd__buf_2
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23518_ _23514_/CLK _23518_/D VGND VGND VPWR VPWR _17684_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24498_ _24042_/CLK _24498_/D HRESETn VGND VGND VPWR VPWR _24498_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ _13955_/Y _14249_/X _14232_/X _14249_/X VGND VGND VPWR VPWR _14251_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17648__A _21336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23449_ _23425_/CLK _19116_/X VGND VGND VPWR VPWR _23449_/Q sky130_fd_sc_hd__dfxtp_4
X_13202_ _13202_/A _18702_/A VGND VGND VPWR VPWR _13202_/X sky130_fd_sc_hd__or2_4
X_14182_ _24829_/Q _14171_/X _24828_/Q _14176_/X VGND VGND VPWR VPWR _14182_/X sky130_fd_sc_hd__o22a_4
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13133_ _13207_/A _13133_/B _13133_/C VGND VGND VPWR VPWR _13133_/X sky130_fd_sc_hd__or3_4
XANTENNA__15168__A _14941_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11696__A _11708_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25119_ _25123_/CLK _12247_/X HRESETn VGND VGND VPWR VPWR _25119_/Q sky130_fd_sc_hd__dfrtp_4
X_18990_ _18990_/A VGND VGND VPWR VPWR _18990_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13064_ _13238_/A _13061_/X _13064_/C VGND VGND VPWR VPWR _13073_/B sky130_fd_sc_hd__and3_4
X_17941_ _17877_/A _23447_/Q VGND VGND VPWR VPWR _17943_/B sky130_fd_sc_hd__or2_4
XANTENNA__21578__A1 _21570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20802__A _20759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12015_ _23796_/Q _12015_/B VGND VGND VPWR VPWR _12016_/B sky130_fd_sc_hd__and2_4
X_17872_ _17968_/A _17872_/B _17872_/C VGND VGND VPWR VPWR _17872_/X sky130_fd_sc_hd__and3_4
XFILLER_26_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23968__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19611_ _19609_/Y _19604_/X _19610_/X _19604_/X VGND VGND VPWR VPWR _19611_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_41_0_HCLK clkbuf_7_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_83_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16823_ _24075_/Q VGND VGND VPWR VPWR _16823_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19542_ _21608_/B _19539_/X _11848_/X _19539_/X VGND VGND VPWR VPWR _19542_/X sky130_fd_sc_hd__a2bb2o_4
X_13966_ _24891_/Q _13944_/B _24891_/Q _13944_/B VGND VGND VPWR VPWR _13967_/A sky130_fd_sc_hd__a2bb2o_4
X_16754_ _15892_/A _16831_/D _15839_/Y _24086_/Q VGND VGND VPWR VPWR _16756_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16206__B1 _15897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12917_ _12802_/Y _12917_/B VGND VGND VPWR VPWR _12920_/B sky130_fd_sc_hd__or2_4
X_15705_ _15693_/X _15689_/X _15704_/X _21567_/A _15661_/A VGND VGND VPWR VPWR _24471_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_19_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16685_ _16685_/A VGND VGND VPWR VPWR _16685_/Y sky130_fd_sc_hd__inv_2
X_19473_ _19467_/Y VGND VGND VPWR VPWR _19473_/X sky130_fd_sc_hd__buf_2
X_13897_ _13854_/X _13897_/B VGND VGND VPWR VPWR _13898_/B sky130_fd_sc_hd__or2_4
XFILLER_62_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18424_ _18422_/Y _18552_/A _18551_/A _18424_/D VGND VGND VPWR VPWR _18427_/C sky130_fd_sc_hd__or4_4
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12848_ _12878_/A VGND VGND VPWR VPWR _12972_/A sky130_fd_sc_hd__buf_2
X_15636_ _15619_/X _15617_/X _15635_/X _20822_/A _15585_/A VGND VGND VPWR VPWR _24502_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_15_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15567_ _15565_/Y _15558_/X _15566_/X _15558_/A VGND VGND VPWR VPWR _15567_/X sky130_fd_sc_hd__a2bb2o_4
X_18355_ _23813_/Q VGND VGND VPWR VPWR _18355_/X sky130_fd_sc_hd__buf_2
X_12779_ _22900_/A VGND VGND VPWR VPWR _12779_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18942__A _17685_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14518_ _14506_/X _14504_/Y _14517_/X _21751_/A _14507_/Y VGND VGND VPWR VPWR _14518_/X
+ sky130_fd_sc_hd__a32o_4
X_17306_ _17306_/A VGND VGND VPWR VPWR _17306_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24756__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15498_ _15482_/X _15483_/X _15497_/X _24560_/Q _15495_/X VGND VGND VPWR VPWR _24560_/D
+ sky130_fd_sc_hd__a32o_4
X_18286_ _23860_/Q _18286_/B VGND VGND VPWR VPWR _18286_/X sky130_fd_sc_hd__or2_4
X_14449_ _21012_/A VGND VGND VPWR VPWR _21008_/A sky130_fd_sc_hd__buf_2
X_17237_ _17237_/A VGND VGND VPWR VPWR _17237_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12990__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19678__A1_N _19677_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17168_ _17031_/A _16858_/A VGND VGND VPWR VPWR _17168_/X sky130_fd_sc_hd__or2_4
XANTENNA__22614__D _22613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16119_ _24327_/Q VGND VGND VPWR VPWR _16119_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16288__A3 _15704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17099_ _24048_/Q _17099_/B VGND VGND VPWR VPWR _17101_/B sky130_fd_sc_hd__or2_4
XFILLER_9_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19809_ _19801_/A _18067_/A _19808_/X _23201_/Q _19802_/A VGND VGND VPWR VPWR _23201_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23638__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22820_ _22820_/A _22638_/X VGND VGND VPWR VPWR _22820_/X sky130_fd_sc_hd__or2_4
XFILLER_42_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_218_0_HCLK clkbuf_8_219_0_HCLK/A VGND VGND VPWR VPWR _24101_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21543__A _21543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13045__B _23076_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22751_ _24245_/Q _21553_/X _20780_/X _22750_/X VGND VGND VPWR VPWR _22751_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21741__B2 _21088_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21702_ _21698_/Y _21699_/X _21700_/X _21701_/X VGND VGND VPWR VPWR _21703_/B sky130_fd_sc_hd__a211o_4
XANTENNA__15541__A _19442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21262__B _21128_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22682_ _16505_/Y _22011_/A _15352_/Y _22452_/X VGND VGND VPWR VPWR _22682_/X sky130_fd_sc_hd__o22a_4
XFILLER_90_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24421_ _24590_/CLK _15843_/X HRESETn VGND VGND VPWR VPWR _24421_/Q sky130_fd_sc_hd__dfrtp_4
X_21633_ _18043_/A _21631_/X _21632_/X VGND VGND VPWR VPWR _21633_/X sky130_fd_sc_hd__and3_4
XANTENNA__24812__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24497__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24352_ _24333_/CLK _24352_/D HRESETn VGND VGND VPWR VPWR _16054_/A sky130_fd_sc_hd__dfrtp_4
X_21564_ _21564_/A _21564_/B VGND VGND VPWR VPWR _21602_/A sky130_fd_sc_hd__nor2_4
XANTENNA__11993__B1 _11607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24426__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23303_ _23303_/CLK _19528_/X VGND VGND VPWR VPWR _23303_/Q sky130_fd_sc_hd__dfxtp_4
X_20515_ _20465_/A VGND VGND VPWR VPWR _20515_/X sky130_fd_sc_hd__buf_2
XANTENNA__15184__B1 _15126_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24283_ _24262_/CLK _24283_/D HRESETn VGND VGND VPWR VPWR _14956_/A sky130_fd_sc_hd__dfrtp_4
X_21495_ _22148_/A _21494_/X VGND VGND VPWR VPWR _21495_/X sky130_fd_sc_hd__or2_4
X_23234_ _23112_/CLK _19725_/X VGND VGND VPWR VPWR _19723_/A sky130_fd_sc_hd__dfxtp_4
X_20446_ _20425_/A VGND VGND VPWR VPWR _20446_/X sky130_fd_sc_hd__buf_2
XFILLER_119_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23165_ _23156_/CLK _23165_/D VGND VGND VPWR VPWR _19908_/A sky130_fd_sc_hd__dfxtp_4
X_20377_ _23674_/Q _20374_/A VGND VGND VPWR VPWR _20377_/Y sky130_fd_sc_hd__nand2_4
XFILLER_106_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22116_ _20753_/A VGND VGND VPWR VPWR _22116_/X sky130_fd_sc_hd__buf_2
XFILLER_133_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23096_ _23249_/CLK _23096_/D VGND VGND VPWR VPWR _20088_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__20622__A _13537_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22047_ _22047_/A _21638_/X VGND VGND VPWR VPWR _22047_/X sky130_fd_sc_hd__or2_4
XFILLER_0_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14977__D _14990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_28_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_28_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25214__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13820_ _13852_/A _13830_/C _13815_/X _13851_/B VGND VGND VPWR VPWR _13820_/X sky130_fd_sc_hd__or4_4
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23998_ _25217_/CLK _17379_/Y HRESETn VGND VGND VPWR VPWR _23998_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13751_ _13717_/B VGND VGND VPWR VPWR _13776_/C sky130_fd_sc_hd__buf_2
X_22949_ _16312_/Y _21896_/X _16050_/Y _22549_/X VGND VGND VPWR VPWR _22949_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13670__B1 _13632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12702_ _12704_/B VGND VGND VPWR VPWR _12703_/B sky130_fd_sc_hd__inv_2
X_16470_ _16469_/Y _16465_/X _16291_/X _16465_/X VGND VGND VPWR VPWR _16470_/X sky130_fd_sc_hd__a2bb2o_4
X_13682_ _23687_/Q VGND VGND VPWR VPWR _13682_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15421_ _16228_/A VGND VGND VPWR VPWR _15421_/X sky130_fd_sc_hd__buf_2
X_12633_ _12591_/X _12632_/X VGND VGND VPWR VPWR _12933_/C sky130_fd_sc_hd__or2_4
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24619_ _24620_/CLK _15307_/X HRESETn VGND VGND VPWR VPWR _24619_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20299__A1 _14223_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15352_ _15352_/A VGND VGND VPWR VPWR _15352_/Y sky130_fd_sc_hd__inv_2
X_18140_ _16102_/A _18213_/D _16058_/Y _23871_/Q VGND VGND VPWR VPWR _18145_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12564_ _12555_/X _12558_/X _12561_/X _12563_/X VGND VGND VPWR VPWR _12591_/B sky130_fd_sc_hd__or4_4
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14303_ HWDATA[1] VGND VGND VPWR VPWR _16216_/A sky130_fd_sc_hd__buf_2
XANTENNA__11984__B1 _11643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11515_ _11514_/X VGND VGND VPWR VPWR _11516_/B sky130_fd_sc_hd__buf_2
X_18071_ _18968_/A _18067_/X _19467_/A VGND VGND VPWR VPWR _18071_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__24167__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15283_ _15281_/Y _15276_/X _15282_/X _15276_/X VGND VGND VPWR VPWR _15283_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12495_ _12495_/A _12495_/B VGND VGND VPWR VPWR _12495_/X sky130_fd_sc_hd__or2_4
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17022_ _17022_/A _17022_/B VGND VGND VPWR VPWR _17055_/A sky130_fd_sc_hd__or2_4
X_14234_ _14234_/A VGND VGND VPWR VPWR _14234_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14165_ _14160_/B _14165_/B VGND VGND VPWR VPWR _14170_/B sky130_fd_sc_hd__or2_4
XFILLER_113_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15478__A1 _15368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22731__B _22952_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13116_ _13054_/X VGND VGND VPWR VPWR _13116_/X sky130_fd_sc_hd__buf_2
XFILLER_112_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14096_ _14096_/A VGND VGND VPWR VPWR _14096_/Y sky130_fd_sc_hd__inv_2
X_18973_ _18972_/Y _18970_/X _18880_/X _18970_/X VGND VGND VPWR VPWR _23501_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16660__A1_N _16658_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13047_ _13047_/A _13045_/X _13047_/C VGND VGND VPWR VPWR _13047_/X sky130_fd_sc_hd__and3_4
X_17924_ _17924_/A _17924_/B VGND VGND VPWR VPWR _17924_/X sky130_fd_sc_hd__or2_4
XANTENNA__16427__B1 _16261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21420__B1 _22351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17855_ _17781_/A _17855_/B VGND VGND VPWR VPWR _17857_/B sky130_fd_sc_hd__or2_4
XFILLER_93_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23731__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16806_ _15830_/Y _24089_/Q _15830_/Y _24089_/Q VGND VGND VPWR VPWR _16806_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17786_ _17727_/A VGND VGND VPWR VPWR _17924_/A sky130_fd_sc_hd__buf_2
XFILLER_54_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14998_ _14881_/A _14995_/X VGND VGND VPWR VPWR _14998_/X sky130_fd_sc_hd__or2_4
XFILLER_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19525_ _23304_/Q VGND VGND VPWR VPWR _19525_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21363__A _21363_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16737_ _23964_/Q VGND VGND VPWR VPWR _17502_/B sky130_fd_sc_hd__inv_2
XFILLER_34_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13949_ _13998_/B VGND VGND VPWR VPWR _13950_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_191_0_HCLK clkbuf_7_95_0_HCLK/X VGND VGND VPWR VPWR _25091_/CLK sky130_fd_sc_hd__clkbuf_1
X_19456_ _21501_/B _19449_/X _19455_/X _19449_/X VGND VGND VPWR VPWR _23330_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21082__B _21082_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24937__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16668_ _14755_/Y _16666_/X _16376_/X _16666_/X VGND VGND VPWR VPWR _24098_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18407_ _18386_/X _18407_/B _18401_/X _18406_/X VGND VGND VPWR VPWR _18408_/B sky130_fd_sc_hd__or4_4
Xclkbuf_8_48_0_HCLK clkbuf_7_24_0_HCLK/X VGND VGND VPWR VPWR _23979_/CLK sky130_fd_sc_hd__clkbuf_1
X_15619_ _16624_/A VGND VGND VPWR VPWR _15619_/X sky130_fd_sc_hd__buf_2
X_19387_ _11635_/A VGND VGND VPWR VPWR _19387_/X sky130_fd_sc_hd__buf_2
X_16599_ _14827_/Y _16595_/X _15501_/X _16595_/X VGND VGND VPWR VPWR _16599_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_5_29_0_HCLK_A clkbuf_4_14_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22906__B _22887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21487__B1 _21172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24590__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18338_ _18420_/A VGND VGND VPWR VPWR _18338_/X sky130_fd_sc_hd__buf_2
XFILLER_124_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15166__B1 _15126_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18269_ _18284_/A _18267_/X _18269_/C VGND VGND VPWR VPWR _23866_/D sky130_fd_sc_hd__and3_4
XFILLER_30_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16613__A1_N _14835_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20300_ _20300_/A VGND VGND VPWR VPWR _23634_/D sky130_fd_sc_hd__inv_2
X_21280_ _21280_/A VGND VGND VPWR VPWR _21280_/X sky130_fd_sc_hd__buf_2
X_20231_ _23773_/Q _20225_/B VGND VGND VPWR VPWR _20257_/B sky130_fd_sc_hd__and2_4
XANTENNA__19852__B1 _19828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15469__A1 _15368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20162_ _23777_/Q _20162_/B VGND VGND VPWR VPWR _20162_/X sky130_fd_sc_hd__or2_4
XFILLER_115_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23819__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16130__A2 _16135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15536__A _15535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20093_ _23094_/Q VGND VGND VPWR VPWR _20093_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24970_ _24750_/CLK _24970_/D HRESETn VGND VGND VPWR VPWR _21696_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_97_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23921_ _24957_/CLK _23921_/D HRESETn VGND VGND VPWR VPWR _11665_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_58_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23852_ _23852_/CLK _18317_/X HRESETn VGND VGND VPWR VPWR _18152_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22803_ _24280_/Q _22616_/X _22351_/X VGND VGND VPWR VPWR _22803_/X sky130_fd_sc_hd__o21a_4
X_23783_ _24980_/CLK _20686_/Y HRESETn VGND VGND VPWR VPWR _11881_/A sky130_fd_sc_hd__dfrtp_4
X_20995_ _21006_/A _19943_/Y VGND VGND VPWR VPWR _20996_/C sky130_fd_sc_hd__or2_4
XFILLER_26_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22911__B1 _25218_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15271__A _15271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24678__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22734_ _22677_/A _22734_/B _22734_/C VGND VGND VPWR VPWR _22734_/X sky130_fd_sc_hd__and3_4
XFILLER_77_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24607__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22665_ _22943_/A _22664_/X VGND VGND VPWR VPWR _22665_/Y sky130_fd_sc_hd__nor2_4
XFILLER_16_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24404_ _24590_/CLK _24404_/D HRESETn VGND VGND VPWR VPWR _24404_/Q sky130_fd_sc_hd__dfrtp_4
X_21616_ _17646_/A VGND VGND VPWR VPWR _21617_/A sky130_fd_sc_hd__buf_2
XFILLER_16_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21720__B _21720_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22596_ _22364_/X _22595_/X _21981_/X _12588_/A _22366_/X VGND VGND VPWR VPWR _22596_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24260__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17203__A2_N _17198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24335_ _24222_/CLK _16101_/X HRESETn VGND VGND VPWR VPWR _24335_/Q sky130_fd_sc_hd__dfrtp_4
X_21547_ _15630_/Y _11986_/X _15797_/Y _21544_/X VGND VGND VPWR VPWR _21547_/X sky130_fd_sc_hd__o22a_4
X_12280_ _12261_/A _12280_/B _12279_/Y VGND VGND VPWR VPWR _25110_/D sky130_fd_sc_hd__and3_4
X_24266_ _24140_/CLK _24266_/D HRESETn VGND VGND VPWR VPWR _22312_/A sky130_fd_sc_hd__dfrtp_4
X_21478_ _21159_/A _19656_/Y VGND VGND VPWR VPWR _21478_/X sky130_fd_sc_hd__or2_4
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23217_ _23401_/CLK _19773_/X VGND VGND VPWR VPWR _23217_/Q sky130_fd_sc_hd__dfxtp_4
X_20429_ _23698_/Q VGND VGND VPWR VPWR _20429_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22442__A2 _20833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24197_ _24197_/CLK _16458_/X HRESETn VGND VGND VPWR VPWR _16457_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16657__B1 _24105_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23148_ _23596_/CLK _19954_/X VGND VGND VPWR VPWR _23148_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_49_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15970_ _15970_/A VGND VGND VPWR VPWR _15970_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23033__A2_N _14428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23079_ _23109_/CLK _23079_/D VGND VGND VPWR VPWR _20127_/A sky130_fd_sc_hd__dfxtp_4
X_14921_ _24679_/Q _24284_/Q _15132_/A _14920_/Y VGND VGND VPWR VPWR _14931_/A sky130_fd_sc_hd__o22a_4
XFILLER_88_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17640_ _17639_/X _17630_/B _17632_/Y VGND VGND VPWR VPWR _17640_/Y sky130_fd_sc_hd__o21ai_4
X_14852_ _14759_/Y VGND VGND VPWR VPWR _15042_/A sky130_fd_sc_hd__buf_2
XANTENNA__15632__A1 _15619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22279__A _22279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15632__B2 _15585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13803_ _13863_/A VGND VGND VPWR VPWR _20164_/A sky130_fd_sc_hd__buf_2
XFILLER_17_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14783_ _24704_/Q _14781_/Y _15022_/A _24113_/Q VGND VGND VPWR VPWR _14784_/D sky130_fd_sc_hd__a2bb2o_4
X_17571_ _17570_/X VGND VGND VPWR VPWR _17572_/B sky130_fd_sc_hd__inv_2
X_11995_ _11990_/A VGND VGND VPWR VPWR _11995_/X sky130_fd_sc_hd__buf_2
XANTENNA__22902__B1 _22564_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19310_ _13141_/B VGND VGND VPWR VPWR _19310_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_201_0_HCLK clkbuf_8_201_0_HCLK/A VGND VGND VPWR VPWR _24596_/CLK sky130_fd_sc_hd__clkbuf_1
X_13734_ _13734_/A VGND VGND VPWR VPWR _13734_/Y sky130_fd_sc_hd__inv_2
X_16522_ _16522_/A VGND VGND VPWR VPWR _16522_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_7_0_HCLK clkbuf_8_7_0_HCLK/A VGND VGND VPWR VPWR _23353_/CLK sky130_fd_sc_hd__clkbuf_1
X_19241_ _19241_/A VGND VGND VPWR VPWR _21927_/B sky130_fd_sc_hd__inv_2
XANTENNA__21911__A _20975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24348__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13665_ _13665_/A VGND VGND VPWR VPWR _13665_/X sky130_fd_sc_hd__buf_2
X_16453_ _16450_/Y _16446_/X _16451_/X _16452_/X VGND VGND VPWR VPWR _24199_/D sky130_fd_sc_hd__a2bb2o_4
X_12616_ _12737_/A _15630_/A _25065_/Q _12615_/Y VGND VGND VPWR VPWR _12616_/X sky130_fd_sc_hd__a2bb2o_4
X_15404_ _15403_/Y _15401_/X _14304_/X _15401_/X VGND VGND VPWR VPWR _15404_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16384_ _16383_/Y _16379_/X _16291_/X _16379_/X VGND VGND VPWR VPWR _16384_/X sky130_fd_sc_hd__a2bb2o_4
X_19172_ _23429_/Q VGND VGND VPWR VPWR _19172_/Y sky130_fd_sc_hd__inv_2
X_13596_ _13558_/A _13558_/B VGND VGND VPWR VPWR _13596_/Y sky130_fd_sc_hd__nand2_4
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15335_ _24611_/Q VGND VGND VPWR VPWR _22884_/A sky130_fd_sc_hd__inv_2
X_18123_ _18122_/Y _18118_/X _18124_/A _18118_/X VGND VGND VPWR VPWR _23881_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15148__B1 _15147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12547_ _12547_/A VGND VGND VPWR VPWR _12547_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15266_ _13745_/B _15260_/X _15240_/A _13722_/X _15262_/X VGND VGND VPWR VPWR _24636_/D
+ sky130_fd_sc_hd__a32o_4
X_18054_ _18045_/X _18046_/X _18050_/X _18053_/X VGND VGND VPWR VPWR _18054_/X sky130_fd_sc_hd__or4_4
XFILLER_8_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12478_ _12412_/B _12478_/B VGND VGND VPWR VPWR _12478_/X sky130_fd_sc_hd__or2_4
X_14217_ _24817_/Q VGND VGND VPWR VPWR _20701_/A sky130_fd_sc_hd__inv_2
X_17005_ _16162_/Y _24049_/Q _16193_/A _16966_/Y VGND VGND VPWR VPWR _17005_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17836__A _17732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15197_ _15197_/A _15197_/B VGND VGND VPWR VPWR _15197_/X sky130_fd_sc_hd__or2_4
XANTENNA__23983__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16648__B1 _22502_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14148_ _24839_/Q _12051_/X _14147_/Y VGND VGND VPWR VPWR _14148_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21358__A _15642_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21641__B1 _23914_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23912__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14079_ _14079_/A VGND VGND VPWR VPWR _14079_/X sky130_fd_sc_hd__buf_2
X_18956_ _18955_/Y _18950_/X _18932_/X _18950_/X VGND VGND VPWR VPWR _18956_/X sky130_fd_sc_hd__a2bb2o_4
X_17907_ _15729_/X _17891_/X _17906_/X _23929_/Q _17765_/X VGND VGND VPWR VPWR _17907_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_79_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18887_ _18886_/Y _18884_/X _18817_/X _18884_/X VGND VGND VPWR VPWR _23531_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17838_ _17934_/A _17838_/B VGND VGND VPWR VPWR _17840_/B sky130_fd_sc_hd__or2_4
Xclkbuf_6_11_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__21093__A _14936_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17769_ _17674_/A VGND VGND VPWR VPWR _17879_/A sky130_fd_sc_hd__buf_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19508_ _23310_/Q VGND VGND VPWR VPWR _19508_/Y sky130_fd_sc_hd__inv_2
X_20780_ _20780_/A VGND VGND VPWR VPWR _20780_/X sky130_fd_sc_hd__buf_2
XFILLER_74_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24089__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24700__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19439_ _14540_/X _19883_/B _19509_/C VGND VGND VPWR VPWR _19440_/A sky130_fd_sc_hd__or3_4
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24018__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22450_ _22450_/A _12063_/X VGND VGND VPWR VPWR _22450_/Y sky130_fd_sc_hd__nor2_4
XFILLER_37_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20437__A _20416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21401_ _21250_/X _21399_/X _13446_/Y _21400_/X VGND VGND VPWR VPWR _21401_/X sky130_fd_sc_hd__a2bb2o_4
X_22381_ _22381_/A _22347_/Y _22381_/C _22380_/X VGND VGND VPWR VPWR HRDATA[12] sky130_fd_sc_hd__or4_4
XANTENNA__22825__A2_N _22822_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20683__A1 _20550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24120_ _24113_/CLK _24120_/D HRESETn VGND VGND VPWR VPWR _14714_/A sky130_fd_sc_hd__dfrtp_4
X_21332_ _21469_/A _21332_/B VGND VGND VPWR VPWR _21334_/B sky130_fd_sc_hd__or2_4
XFILLER_135_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20683__B2 _20602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22652__A _21064_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14892__A2_N _24280_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24051_ _24049_/CLK _24051_/D HRESETn VGND VGND VPWR VPWR _24051_/Q sky130_fd_sc_hd__dfrtp_4
X_21263_ _12349_/A _21408_/B VGND VGND VPWR VPWR _21263_/X sky130_fd_sc_hd__or2_4
XFILLER_132_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16650__A _16643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20435__A1 _15395_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23002_ _23002_/A _22834_/B VGND VGND VPWR VPWR _23002_/X sky130_fd_sc_hd__or2_4
X_20214_ _23771_/Q _20225_/B VGND VGND VPWR VPWR _20224_/B sky130_fd_sc_hd__and2_4
XANTENNA__23653__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21194_ _21237_/A VGND VGND VPWR VPWR _21500_/A sky130_fd_sc_hd__buf_2
XFILLER_103_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20145_ _23072_/Q VGND VGND VPWR VPWR _20145_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15311__B1 HADDR[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16654__A3 _11585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24953_ _24953_/CLK _24953_/D HRESETn VGND VGND VPWR VPWR _11657_/A sky130_fd_sc_hd__dfrtp_4
X_20076_ _20076_/A VGND VGND VPWR VPWR _20076_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12402__B _12448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20900__A _20900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17481__A _17481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24859__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23904_ _24928_/CLK _23904_/D HRESETn VGND VGND VPWR VPWR _23904_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24884_ _24884_/CLK _24884_/D HRESETn VGND VGND VPWR VPWR _24884_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12428__A1 _12391_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22397__A1_N _12498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23835_ _23826_/CLK _18483_/Y HRESETn VGND VGND VPWR VPWR _23835_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11780_ _25180_/Q VGND VGND VPWR VPWR _11780_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23766_ _24643_/CLK _20259_/X HRESETn VGND VGND VPWR VPWR _23766_/Q sky130_fd_sc_hd__dfrtp_4
X_20978_ _20978_/A _20978_/B VGND VGND VPWR VPWR _20978_/X sky130_fd_sc_hd__or2_4
XFILLER_54_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24441__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22717_ _22360_/X _22702_/X _22705_/X _22711_/X _22716_/X VGND VGND VPWR VPWR _22718_/D
+ sky130_fd_sc_hd__o41a_4
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15917__A2 _15915_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23697_ _24349_/CLK _20428_/Y HRESETn VGND VGND VPWR VPWR _13498_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_41_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13450_ _24938_/Q VGND VGND VPWR VPWR _13450_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19201__A _18678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_31_0_HCLK clkbuf_8_31_0_HCLK/A VGND VGND VPWR VPWR _23908_/CLK sky130_fd_sc_hd__clkbuf_1
X_22648_ _22129_/X _22645_/X _22646_/X _24414_/Q _22647_/X VGND VGND VPWR VPWR _22648_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20030__A2_N _20027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12401_ _12433_/A _12401_/B VGND VGND VPWR VPWR _12401_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_94_0_HCLK clkbuf_8_95_0_HCLK/A VGND VGND VPWR VPWR _23680_/CLK sky130_fd_sc_hd__clkbuf_1
X_13381_ _24977_/Q VGND VGND VPWR VPWR _13381_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22663__A2 _20910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22579_ _22691_/A _22579_/B _22579_/C VGND VGND VPWR VPWR _22614_/A sky130_fd_sc_hd__and3_4
X_15120_ _24681_/Q _15119_/Y VGND VGND VPWR VPWR _15120_/X sky130_fd_sc_hd__or2_4
X_12332_ _24491_/Q VGND VGND VPWR VPWR _12332_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24318_ _24055_/CLK _16146_/X HRESETn VGND VGND VPWR VPWR _24318_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20674__B2 _20602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22562__A _22677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15051_ _15051_/A VGND VGND VPWR VPWR _15051_/Y sky130_fd_sc_hd__inv_2
X_12263_ _12262_/X VGND VGND VPWR VPWR _12263_/Y sky130_fd_sc_hd__inv_2
X_24249_ _24225_/CLK _24249_/D HRESETn VGND VGND VPWR VPWR _24249_/Q sky130_fd_sc_hd__dfrtp_4
X_14002_ _13996_/Y _13937_/X _13938_/X _14001_/X VGND VGND VPWR VPWR _14002_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21178__A _21178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12194_ _12165_/X VGND VGND VPWR VPWR _12538_/B sky130_fd_sc_hd__inv_2
XANTENNA__19292__B2 _19289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18810_ _18806_/Y _18809_/X _18764_/X _18809_/X VGND VGND VPWR VPWR _18810_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14105__A1 _23126_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15302__B1 HWRITE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19790_ _23210_/Q VGND VGND VPWR VPWR _21522_/B sky130_fd_sc_hd__inv_2
XANTENNA__17094__C _17132_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22179__A1 _12098_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22179__B2 _22228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18741_ _18738_/Y _18736_/X _18740_/X _18736_/X VGND VGND VPWR VPWR _23581_/D sky130_fd_sc_hd__a2bb2o_4
X_15953_ _15928_/X VGND VGND VPWR VPWR _15953_/X sky130_fd_sc_hd__buf_2
X_14904_ _14903_/Y _24255_/Q _14903_/Y _24255_/Q VGND VGND VPWR VPWR _14904_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15904__A _24397_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18672_ _23604_/Q VGND VGND VPWR VPWR _18672_/Y sky130_fd_sc_hd__inv_2
X_15884_ _24404_/Q VGND VGND VPWR VPWR _15884_/Y sky130_fd_sc_hd__inv_2
X_17623_ _17619_/A _17614_/B _17622_/X VGND VGND VPWR VPWR _23942_/D sky130_fd_sc_hd__and3_4
XFILLER_56_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24529__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14835_ _24129_/Q VGND VGND VPWR VPWR _14835_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17554_ _16692_/Y _17554_/B VGND VGND VPWR VPWR _17554_/X sky130_fd_sc_hd__or2_4
X_11978_ _11965_/Y VGND VGND VPWR VPWR _11978_/X sky130_fd_sc_hd__buf_2
X_14766_ _14765_/Y VGND VGND VPWR VPWR _15004_/A sky130_fd_sc_hd__buf_2
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16505_ _16505_/A VGND VGND VPWR VPWR _16505_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24182__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13717_ _13753_/A _13717_/B _13716_/X VGND VGND VPWR VPWR _13766_/D sky130_fd_sc_hd__or3_4
X_14697_ _24713_/Q VGND VGND VPWR VPWR _14697_/Y sky130_fd_sc_hd__inv_2
X_17485_ _22307_/A VGND VGND VPWR VPWR _17486_/A sky130_fd_sc_hd__inv_2
X_19224_ _19223_/Y _19218_/X _19201_/X _19218_/X VGND VGND VPWR VPWR _23410_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22918__A1_N _21546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24111__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16436_ _24205_/Q VGND VGND VPWR VPWR _16436_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13648_ _13647_/Y VGND VGND VPWR VPWR _13649_/A sky130_fd_sc_hd__buf_2
XFILLER_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19155_ _19155_/A VGND VGND VPWR VPWR _19155_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13579_ _13571_/X _13553_/X _13578_/X _13576_/X _11653_/A VGND VGND VPWR VPWR _24959_/D
+ sky130_fd_sc_hd__a32o_4
X_16367_ _16366_/Y _16364_/X _15982_/X _16364_/X VGND VGND VPWR VPWR _24230_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_2_0_HCLK clkbuf_5_2_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_18106_ _18093_/A _18092_/X VGND VGND VPWR VPWR _18106_/X sky130_fd_sc_hd__or2_4
X_15318_ _16231_/A _20926_/A VGND VGND VPWR VPWR _15531_/B sky130_fd_sc_hd__or2_4
XFILLER_34_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16298_ _18263_/A VGND VGND VPWR VPWR _18258_/A sky130_fd_sc_hd__buf_2
X_19086_ _17828_/B VGND VGND VPWR VPWR _19086_/Y sky130_fd_sc_hd__inv_2
X_18037_ _17625_/A _18036_/X _18025_/D _18061_/B VGND VGND VPWR VPWR _23902_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17566__A _16718_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15249_ _14099_/A VGND VGND VPWR VPWR _15250_/A sky130_fd_sc_hd__buf_2
XANTENNA__12355__B1 _12403_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16097__B2 _16090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19988_ _23134_/Q VGND VGND VPWR VPWR _19988_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18939_ _18937_/Y _18935_/X _18938_/X _18935_/X VGND VGND VPWR VPWR _23512_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21816__A _20966_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21950_ _21211_/A _21950_/B VGND VGND VPWR VPWR _21950_/X sky130_fd_sc_hd__or2_4
XFILLER_55_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24952__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20901_ _22587_/B VGND VGND VPWR VPWR _22497_/B sky130_fd_sc_hd__buf_2
X_21881_ _21881_/A VGND VGND VPWR VPWR _21881_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13334__A _20818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23620_ _24897_/CLK _23620_/D HRESETn VGND VGND VPWR VPWR _20175_/A sky130_fd_sc_hd__dfrtp_4
X_20832_ _20832_/A VGND VGND VPWR VPWR _22858_/A sky130_fd_sc_hd__buf_2
XFILLER_54_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22647__A _22992_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22342__B2 _21870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18010__A2 _15915_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23551_ _24998_/CLK _18829_/X VGND VGND VPWR VPWR _18827_/A sky130_fd_sc_hd__dfxtp_4
X_20763_ _11940_/Y VGND VGND VPWR VPWR _21591_/B sky130_fd_sc_hd__buf_2
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22502_ _22502_/A _22580_/B VGND VGND VPWR VPWR _22502_/X sky130_fd_sc_hd__or2_4
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_18_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23482_ _23482_/CLK _23482_/D VGND VGND VPWR VPWR _23482_/Q sky130_fd_sc_hd__dfxtp_4
X_20694_ _12022_/A _20695_/B VGND VGND VPWR VPWR _20694_/X sky130_fd_sc_hd__and2_4
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25221_ _24405_/CLK _23043_/X HRESETn VGND VGND VPWR VPWR _25221_/Q sky130_fd_sc_hd__dfrtp_4
X_22433_ _22433_/A _22433_/B _22432_/X VGND VGND VPWR VPWR _22457_/C sky130_fd_sc_hd__and3_4
XFILLER_17_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21853__B1 _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25152_ _24824_/CLK _25152_/D HRESETn VGND VGND VPWR VPWR _25152_/Q sky130_fd_sc_hd__dfrtp_4
X_22364_ _20753_/A VGND VGND VPWR VPWR _22364_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23834__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20120__A3 _13665_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25058__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24103_ _24138_/CLK _16661_/X HRESETn VGND VGND VPWR VPWR _14709_/A sky130_fd_sc_hd__dfrtp_4
X_21315_ _14036_/Y _14015_/A _14059_/A _20844_/B VGND VGND VPWR VPWR _21315_/X sky130_fd_sc_hd__a2bb2o_4
X_25083_ _25091_/CLK _12499_/X HRESETn VGND VGND VPWR VPWR _12497_/A sky130_fd_sc_hd__dfrtp_4
X_22295_ _20909_/X _22294_/X _22240_/X _25201_/Q _21402_/X VGND VGND VPWR VPWR _22295_/X
+ sky130_fd_sc_hd__a32o_4
X_24034_ _24031_/CLK _24034_/D HRESETn VGND VGND VPWR VPWR _24034_/Q sky130_fd_sc_hd__dfrtp_4
X_21246_ _21245_/X VGND VGND VPWR VPWR _21246_/X sky130_fd_sc_hd__buf_2
XFILLER_117_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17285__B1 _25218_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13509__A _13509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21177_ _20753_/A VGND VGND VPWR VPWR _21178_/A sky130_fd_sc_hd__buf_2
XFILLER_133_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20128_ _20127_/Y _20123_/Y _19963_/X _20123_/Y VGND VGND VPWR VPWR _23079_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12950_ _12947_/B VGND VGND VPWR VPWR _12951_/B sky130_fd_sc_hd__inv_2
XANTENNA__24693__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20059_ _20055_/X VGND VGND VPWR VPWR _20060_/A sky130_fd_sc_hd__inv_2
X_24936_ _24937_/CLK _13656_/X HRESETn VGND VGND VPWR VPWR _13655_/A sky130_fd_sc_hd__dfrtp_4
X_11901_ _13368_/A _11900_/Y _13368_/A _11900_/Y VGND VGND VPWR VPWR _11901_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24622__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12881_ _12796_/Y _12947_/A _12809_/Y _12785_/A VGND VGND VPWR VPWR _12881_/X sky130_fd_sc_hd__or4_4
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20592__B1 _20583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24867_ _24870_/CLK _14058_/X HRESETn VGND VGND VPWR VPWR _24867_/Q sky130_fd_sc_hd__dfstp_4
X_11832_ _11827_/Y _11831_/X RsRx_S1 _11831_/X VGND VGND VPWR VPWR _25176_/D sky130_fd_sc_hd__a2bb2o_4
X_14620_ _14620_/A VGND VGND VPWR VPWR _14620_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23818_ _23824_/CLK _23818_/D HRESETn VGND VGND VPWR VPWR _23818_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14271__B1 _14232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24798_ _24859_/CLK _24798_/D HRESETn VGND VGND VPWR VPWR _14270_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_14_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22557__A _22992_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18537__B1 _18449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14452_/X _14437_/X _14549_/X VGND VGND VPWR VPWR _24739_/D sky130_fd_sc_hd__o21a_4
XPHY_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11763_/A _18065_/B _11763_/C _11763_/D VGND VGND VPWR VPWR _11763_/X sky130_fd_sc_hd__or4_4
XFILLER_109_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23749_ _24180_/CLK _23749_/D HRESETn VGND VGND VPWR VPWR _23749_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _23698_/Q _13501_/Y VGND VGND VPWR VPWR _13503_/B sky130_fd_sc_hd__or2_4
XFILLER_41_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14482_/A VGND VGND VPWR VPWR _14482_/X sky130_fd_sc_hd__buf_2
X_17270_ _17270_/A VGND VGND VPWR VPWR _17270_/Y sky130_fd_sc_hd__inv_2
XPHY_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11660_/X _11669_/X _11694_/C _11694_/D VGND VGND VPWR VPWR _11694_/X sky130_fd_sc_hd__or4_4
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15220__C1 _15147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13433_ _24935_/Q _13432_/A _22271_/A _13432_/Y VGND VGND VPWR VPWR _13440_/B sky130_fd_sc_hd__o22a_4
X_16221_ _14369_/B _14435_/D _16221_/C VGND VGND VPWR VPWR _16221_/X sky130_fd_sc_hd__and3_4
XPHY_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15771__B1 _15770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16152_ _16165_/A VGND VGND VPWR VPWR _16152_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13364_ _11913_/Y _13363_/X _11604_/X _13363_/X VGND VGND VPWR VPWR _13364_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12315_ _12474_/C _24483_/Q _12412_/D _24483_/Q VGND VGND VPWR VPWR _12315_/X sky130_fd_sc_hd__a2bb2o_4
X_15103_ _14946_/Y _15136_/C VGND VGND VPWR VPWR _15103_/X sky130_fd_sc_hd__or2_4
X_16083_ _16083_/A VGND VGND VPWR VPWR _16084_/A sky130_fd_sc_hd__buf_2
XANTENNA__17386__A _17270_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15523__B1 _24548_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13295_ _13159_/X _13293_/X _13295_/C VGND VGND VPWR VPWR _13296_/C sky130_fd_sc_hd__and3_4
XANTENNA__16290__A HWDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15034_ _15034_/A _15034_/B VGND VGND VPWR VPWR _15034_/X sky130_fd_sc_hd__or2_4
X_19911_ _19918_/A VGND VGND VPWR VPWR _19911_/X sky130_fd_sc_hd__buf_2
X_12246_ _12174_/B _12243_/B VGND VGND VPWR VPWR _12246_/Y sky130_fd_sc_hd__nand2_4
XFILLER_123_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19804__A3 _13665_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19842_ _19841_/X VGND VGND VPWR VPWR _19842_/X sky130_fd_sc_hd__buf_2
X_12177_ _12177_/A VGND VGND VPWR VPWR _12275_/A sky130_fd_sc_hd__inv_2
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21636__A _20745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19773_ _21329_/B _19772_/X _19728_/X _19772_/X VGND VGND VPWR VPWR _19773_/X sky130_fd_sc_hd__a2bb2o_4
X_16985_ _24318_/Q _24056_/Q _16143_/Y _17022_/A VGND VGND VPWR VPWR _16990_/B sky130_fd_sc_hd__o22a_4
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18724_ _18719_/A VGND VGND VPWR VPWR _18724_/X sky130_fd_sc_hd__buf_2
XFILLER_114_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22021__B1 _22497_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15936_ _15928_/X VGND VGND VPWR VPWR _15936_/X sky130_fd_sc_hd__buf_2
XFILLER_76_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24363__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18655_ _21508_/B _18650_/X _15559_/X _18650_/X VGND VGND VPWR VPWR _18655_/X sky130_fd_sc_hd__a2bb2o_4
X_15867_ _15826_/A VGND VGND VPWR VPWR _15885_/A sky130_fd_sc_hd__buf_2
XFILLER_97_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17606_ _16685_/Y _17594_/B VGND VGND VPWR VPWR _17606_/Y sky130_fd_sc_hd__nand2_4
X_14818_ _14818_/A VGND VGND VPWR VPWR _14818_/Y sky130_fd_sc_hd__inv_2
X_18586_ _24239_/Q _18495_/B _16361_/Y _23823_/Q VGND VGND VPWR VPWR _18587_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15798_ _15797_/Y _15795_/X _15279_/X _15795_/X VGND VGND VPWR VPWR _24433_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17537_ _17483_/A _17535_/A VGND VGND VPWR VPWR _17537_/X sky130_fd_sc_hd__or2_4
X_14749_ _14749_/A _14749_/B _14745_/X _14748_/X VGND VGND VPWR VPWR _14749_/X sky130_fd_sc_hd__or4_4
XANTENNA__16465__A _16401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18595__A1_N _16351_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17200__B1 _17199_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17468_ _17468_/A VGND VGND VPWR VPWR _17468_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19207_ _18801_/X VGND VGND VPWR VPWR _19207_/X sky130_fd_sc_hd__buf_2
X_16419_ _16418_/Y _16414_/X _16254_/X _16414_/X VGND VGND VPWR VPWR _16419_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15762__B1 _15761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17399_ _17329_/A _17325_/C VGND VGND VPWR VPWR _17399_/X sky130_fd_sc_hd__or2_4
X_19138_ _19136_/Y _19137_/X _19115_/X _19137_/X VGND VGND VPWR VPWR _19138_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25151__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19069_ _19068_/Y _19064_/X _18932_/X _19064_/X VGND VGND VPWR VPWR _23466_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15606__A1_N _12617_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14713__A _24114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21100_ _14754_/Y _22017_/A VGND VGND VPWR VPWR _21100_/X sky130_fd_sc_hd__or2_4
XFILLER_133_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22080_ _21519_/A _22078_/X _22079_/X VGND VGND VPWR VPWR _22080_/X sky130_fd_sc_hd__and3_4
XANTENNA__17446__D _11720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21031_ _20786_/A VGND VGND VPWR VPWR _21408_/B sky130_fd_sc_hd__buf_2
XANTENNA__13329__A _15422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15544__A _19448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22982_ _22982_/A _22982_/B _22980_/X _22982_/D VGND VGND VPWR VPWR _22982_/X sky130_fd_sc_hd__or4_4
XFILLER_41_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18767__B1 _18740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21933_ _20980_/A _21933_/B _21932_/X VGND VGND VPWR VPWR _21933_/X sky130_fd_sc_hd__and3_4
X_24721_ _24723_/CLK _14669_/X HRESETn VGND VGND VPWR VPWR _24721_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24033__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24652_ _24654_/CLK _24652_/D HRESETn VGND VGND VPWR VPWR _14925_/A sky130_fd_sc_hd__dfrtp_4
X_21864_ _22279_/A VGND VGND VPWR VPWR _21864_/X sky130_fd_sc_hd__buf_2
XFILLER_15_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22315__B2 _16305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23603_ _24008_/CLK _23603_/D VGND VGND VPWR VPWR _23603_/Q sky130_fd_sc_hd__dfxtp_4
X_20815_ _20814_/X VGND VGND VPWR VPWR _20815_/X sky130_fd_sc_hd__buf_2
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24583_ _24017_/CLK _15419_/X HRESETn VGND VGND VPWR VPWR _20741_/B sky130_fd_sc_hd__dfrtp_4
X_21795_ _21795_/A _21795_/B VGND VGND VPWR VPWR _21795_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__22866__A2 _16134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19192__B1 _19170_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23534_ _23457_/CLK _18878_/X VGND VGND VPWR VPWR _17681_/B sky130_fd_sc_hd__dfxtp_4
X_20746_ _20745_/X VGND VGND VPWR VPWR _22201_/A sky130_fd_sc_hd__buf_2
XFILLER_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23465_ _23419_/CLK _23465_/D VGND VGND VPWR VPWR _17880_/B sky130_fd_sc_hd__dfxtp_4
X_20677_ _20675_/Y _20672_/Y _20676_/X VGND VGND VPWR VPWR _20677_/X sky130_fd_sc_hd__o21a_4
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25204_ _24385_/CLK _25204_/D HRESETn VGND VGND VPWR VPWR _11583_/A sky130_fd_sc_hd__dfrtp_4
X_22416_ _22495_/A _22416_/B _22416_/C _22416_/D VGND VGND VPWR VPWR _22416_/X sky130_fd_sc_hd__or4_4
X_23396_ _23411_/CLK _23396_/D VGND VGND VPWR VPWR _19265_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_105_0_HCLK clkbuf_7_52_0_HCLK/X VGND VGND VPWR VPWR _24399_/CLK sky130_fd_sc_hd__clkbuf_1
X_25135_ _24974_/CLK _25135_/D HRESETn VGND VGND VPWR VPWR _25135_/Q sky130_fd_sc_hd__dfrtp_4
X_22347_ _22346_/X VGND VGND VPWR VPWR _22347_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_168_0_HCLK clkbuf_7_84_0_HCLK/X VGND VGND VPWR VPWR _23332_/CLK sky130_fd_sc_hd__clkbuf_1
X_12100_ _25126_/Q VGND VGND VPWR VPWR _12219_/A sky130_fd_sc_hd__inv_2
X_13080_ _13203_/A _13080_/B _13079_/X VGND VGND VPWR VPWR _13087_/B sky130_fd_sc_hd__and3_4
X_25066_ _25046_/CLK _25066_/D HRESETn VGND VGND VPWR VPWR _25066_/Q sky130_fd_sc_hd__dfrtp_4
X_22278_ _22278_/A _22188_/X VGND VGND VPWR VPWR _22278_/X sky130_fd_sc_hd__and2_4
XANTENNA__19247__B2 _19244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22840__A _22840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19753__A2_N _19750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12031_ _20696_/A VGND VGND VPWR VPWR _12031_/Y sky130_fd_sc_hd__inv_2
X_24017_ _24017_/CLK _24017_/D HRESETn VGND VGND VPWR VPWR _24017_/Q sky130_fd_sc_hd__dfrtp_4
X_21229_ _21229_/A _21229_/B VGND VGND VPWR VPWR _21230_/C sky130_fd_sc_hd__or2_4
XANTENNA__24874__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15808__A1 _16222_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22026__A2_N _12063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18468__C _18468_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16770_ _15846_/A _24083_/Q _15846_/Y _16769_/Y VGND VGND VPWR VPWR _16770_/X sky130_fd_sc_hd__o22a_4
X_13982_ _13973_/X _13981_/Y _14223_/A _13973_/X VGND VGND VPWR VPWR _13982_/X sky130_fd_sc_hd__a2bb2o_4
X_15721_ _15807_/A _15718_/Y _15720_/X _13458_/B VGND VGND VPWR VPWR _15722_/C sky130_fd_sc_hd__a211o_4
XFILLER_74_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12933_ _12836_/Y _12964_/A _12933_/C _12933_/D VGND VGND VPWR VPWR _12955_/B sky130_fd_sc_hd__or4_4
XFILLER_111_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24919_ _24923_/CLK _13699_/X HRESETn VGND VGND VPWR VPWR _21733_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_74_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18440_ _18440_/A _18440_/B _18459_/A _18446_/A VGND VGND VPWR VPWR _18440_/X sky130_fd_sc_hd__or4_4
X_15652_ _13614_/A VGND VGND VPWR VPWR _21092_/B sky130_fd_sc_hd__inv_2
XFILLER_34_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12864_ _12863_/Y _21980_/A _12858_/X _24432_/Q VGND VGND VPWR VPWR _12864_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14244__B1 _14213_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15587__A3 _15468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14603_ _19946_/C _19167_/B _19946_/C _19167_/B VGND VGND VPWR VPWR _14603_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21191__A _11720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11815_ _25180_/Q _11828_/B _11815_/C _11814_/Y VGND VGND VPWR VPWR _11815_/X sky130_fd_sc_hd__or4_4
X_18371_ _24219_/Q _23842_/Q _16400_/Y _18412_/A VGND VGND VPWR VPWR _18371_/X sky130_fd_sc_hd__o22a_4
X_12795_ _12795_/A _12789_/X _12795_/C _12795_/D VGND VGND VPWR VPWR _12822_/B sky130_fd_sc_hd__or4_4
X_15583_ _11986_/X _15741_/B VGND VGND VPWR VPWR _15584_/A sky130_fd_sc_hd__or2_4
XPHY_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _23978_/Q VGND VGND VPWR VPWR _17323_/D sky130_fd_sc_hd__inv_2
XANTENNA__20868__A1 _22444_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _23896_/Q VGND VGND VPWR VPWR _11746_/Y sky130_fd_sc_hd__inv_2
X_14534_ _21009_/A VGND VGND VPWR VPWR _21205_/A sky130_fd_sc_hd__buf_2
XANTENNA__23756__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18930__B1 _18817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14547__A1 _14482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17253_ _17253_/A VGND VGND VPWR VPWR _17413_/A sky130_fd_sc_hd__inv_2
XANTENNA__19596__A _19613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _11677_/A VGND VGND VPWR VPWR _11677_/Y sky130_fd_sc_hd__inv_2
X_14465_ _19779_/B _14446_/X VGND VGND VPWR VPWR _14465_/X sky130_fd_sc_hd__and2_4
XANTENNA__14547__B2 _14437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19706__A2_N _19701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16204_ _16202_/Y _16203_/X _15894_/X _16203_/X VGND VGND VPWR VPWR _24295_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13416_ _13416_/A VGND VGND VPWR VPWR _14385_/A sky130_fd_sc_hd__inv_2
Xclkbuf_7_64_0_HCLK clkbuf_6_32_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_64_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14396_ _14394_/X _14371_/X _14395_/X _13608_/X _14387_/C VGND VGND VPWR VPWR _14396_/X
+ sky130_fd_sc_hd__a32o_4
X_17184_ _17186_/B VGND VGND VPWR VPWR _17184_/Y sky130_fd_sc_hd__inv_2
X_13347_ _13346_/Y _13344_/X _11626_/X _13344_/X VGND VGND VPWR VPWR _13347_/X sky130_fd_sc_hd__a2bb2o_4
X_16135_ _16134_/X _16135_/B VGND VGND VPWR VPWR _16135_/X sky130_fd_sc_hd__and2_4
XFILLER_6_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13278_ _13278_/A _13276_/X _13278_/C VGND VGND VPWR VPWR _13278_/X sky130_fd_sc_hd__and3_4
X_16066_ _24347_/Q VGND VGND VPWR VPWR _16066_/Y sky130_fd_sc_hd__inv_2
X_12229_ _12175_/C _12228_/X VGND VGND VPWR VPWR _12229_/X sky130_fd_sc_hd__or2_4
X_15017_ _15017_/A VGND VGND VPWR VPWR _24704_/D sky130_fd_sc_hd__inv_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22151__A1_N _11680_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21596__A2 _21109_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19825_ _19825_/A VGND VGND VPWR VPWR _19825_/X sky130_fd_sc_hd__buf_2
XANTENNA__22793__B2 _22548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24544__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12988__A _12992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19756_ _20974_/B _19750_/X _19755_/X _19737_/Y VGND VGND VPWR VPWR _23223_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16968_ _24048_/Q VGND VGND VPWR VPWR _16968_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22545__A1 _21529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18707_ _18704_/Y _18705_/X _18706_/X _18705_/X VGND VGND VPWR VPWR _23593_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22545__B2 _22544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15919_ _15655_/A VGND VGND VPWR VPWR _15919_/X sky130_fd_sc_hd__buf_2
XANTENNA__19278__A1_N _21251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19687_ _18018_/X _19282_/B _19531_/X VGND VGND VPWR VPWR _19688_/A sky130_fd_sc_hd__or3_4
X_16899_ _16784_/Y _16902_/B VGND VGND VPWR VPWR _16900_/B sky130_fd_sc_hd__or2_4
X_18638_ _18638_/A _18638_/B _18637_/Y _11719_/B VGND VGND VPWR VPWR _18638_/X sky130_fd_sc_hd__or4_4
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16775__A2 _16774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18569_ _16381_/Y _23816_/Q _16381_/Y _23816_/Q VGND VGND VPWR VPWR _18569_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15983__B1 _15982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14786__B2 _14754_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20600_ _23737_/Q _13534_/B _20599_/Y VGND VGND VPWR VPWR _20600_/Y sky130_fd_sc_hd__a21oi_4
X_21580_ _21580_/A _11499_/A VGND VGND VPWR VPWR _21580_/X sky130_fd_sc_hd__or2_4
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20531_ _13512_/X VGND VGND VPWR VPWR _20531_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23250_ _23242_/CLK _23250_/D VGND VGND VPWR VPWR _19677_/A sky130_fd_sc_hd__dfxtp_4
X_20462_ _20469_/B VGND VGND VPWR VPWR _20462_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22201_ _22201_/A _22201_/B _22190_/X _22200_/X VGND VGND VPWR VPWR _22201_/X sky130_fd_sc_hd__or4_4
XFILLER_101_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23181_ _23179_/CLK _23181_/D VGND VGND VPWR VPWR _23181_/Q sky130_fd_sc_hd__dfxtp_4
X_20393_ _20393_/A _17187_/X VGND VGND VPWR VPWR _20393_/X sky130_fd_sc_hd__or2_4
XFILLER_119_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22132_ _20838_/X _22128_/Y _20815_/X _22131_/X VGND VGND VPWR VPWR _22132_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15502__A3 _15501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22063_ _22055_/X _19438_/Y VGND VGND VPWR VPWR _22063_/X sky130_fd_sc_hd__or2_4
XFILLER_88_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17754__A _17742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22784__A1 _25214_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21014_ _21006_/A _19922_/Y VGND VGND VPWR VPWR _21014_/X sky130_fd_sc_hd__or2_4
XFILLER_102_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24285__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20795__B1 _20782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24214__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20547__B1 _13515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22965_ _22943_/Y _22965_/B _22951_/Y _22964_/X VGND VGND VPWR VPWR HRDATA[29] sky130_fd_sc_hd__or4_4
X_24704_ _24706_/CLK _24704_/D HRESETn VGND VGND VPWR VPWR _24704_/Q sky130_fd_sc_hd__dfrtp_4
X_21916_ _21924_/A _21916_/B VGND VGND VPWR VPWR _21916_/X sky130_fd_sc_hd__or2_4
X_22896_ _22895_/X VGND VGND VPWR VPWR _22896_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21847_ _21565_/A _21847_/B VGND VGND VPWR VPWR _21855_/B sky130_fd_sc_hd__and2_4
X_24635_ _23762_/CLK _24635_/D HRESETn VGND VGND VPWR VPWR _24635_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15974__B1 _11598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ _11596_/Y _11588_/X _11598_/X _11599_/X VGND VGND VPWR VPWR _11600_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _25066_/Q _12579_/A _12578_/Y _12579_/Y VGND VGND VPWR VPWR _12580_/X sky130_fd_sc_hd__o22a_4
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24566_ _24566_/CLK _24566_/D HRESETn VGND VGND VPWR VPWR _12088_/A sky130_fd_sc_hd__dfrtp_4
X_21778_ _21383_/A _21778_/B VGND VGND VPWR VPWR _21779_/C sky130_fd_sc_hd__or2_4
XFILLER_24_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25073__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ _11530_/X VGND VGND VPWR VPWR _11532_/A sky130_fd_sc_hd__buf_2
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20729_ _20729_/A _20729_/B _23666_/Q VGND VGND VPWR VPWR _20729_/X sky130_fd_sc_hd__or3_4
XFILLER_8_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23517_ _23514_/CLK _23517_/D VGND VGND VPWR VPWR _23517_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24497_ _24042_/CLK _24497_/D HRESETn VGND VGND VPWR VPWR _22975_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25002__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ _14247_/Y _14249_/X _14228_/X _14249_/X VGND VGND VPWR VPWR _14250_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23448_ _23440_/CLK _23448_/D VGND VGND VPWR VPWR _23448_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ _13127_/A _23072_/Q VGND VGND VPWR VPWR _13201_/X sky130_fd_sc_hd__or2_4
XFILLER_137_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14181_ _14175_/X _14179_/X _25154_/Q _14180_/X VGND VGND VPWR VPWR _24830_/D sky130_fd_sc_hd__o22a_4
X_23379_ _23374_/CLK _23379_/D VGND VGND VPWR VPWR _13178_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_125_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13132_ _13171_/A _13130_/X _13131_/X VGND VGND VPWR VPWR _13133_/C sky130_fd_sc_hd__and3_4
XFILLER_87_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14769__A1_N _15034_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25118_ _25123_/CLK _25118_/D HRESETn VGND VGND VPWR VPWR _12082_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_87_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13063_ _13202_/A _13063_/B VGND VGND VPWR VPWR _13064_/C sky130_fd_sc_hd__or2_4
X_17940_ _17705_/X _17939_/X _23927_/Q _17767_/A VGND VGND VPWR VPWR _17940_/X sky130_fd_sc_hd__o22a_4
XFILLER_112_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25049_ _25050_/CLK _12734_/Y HRESETn VGND VGND VPWR VPWR _25049_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14701__B2 _14714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12014_ _23795_/Q _12014_/B VGND VGND VPWR VPWR _12015_/B sky130_fd_sc_hd__and2_4
XANTENNA__21186__A _21109_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17871_ _17903_/A _17871_/B VGND VGND VPWR VPWR _17872_/C sky130_fd_sc_hd__or2_4
XFILLER_79_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_6_0_HCLK clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19610_ _19610_/A VGND VGND VPWR VPWR _19610_/X sky130_fd_sc_hd__buf_2
X_16822_ _16822_/A _16802_/Y VGND VGND VPWR VPWR _16822_/X sky130_fd_sc_hd__or2_4
XFILLER_19_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19541_ _23299_/Q VGND VGND VPWR VPWR _21608_/B sky130_fd_sc_hd__inv_2
X_16753_ _24065_/Q VGND VGND VPWR VPWR _16831_/D sky130_fd_sc_hd__inv_2
XANTENNA__21914__A _20980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13965_ _13952_/X _13964_/Y _24892_/Q _13952_/X VGND VGND VPWR VPWR _13965_/X sky130_fd_sc_hd__a2bb2o_4
X_15704_ _11625_/A VGND VGND VPWR VPWR _15704_/X sky130_fd_sc_hd__buf_2
XFILLER_111_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15912__A _15431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12916_ _12838_/Y _12916_/B VGND VGND VPWR VPWR _12917_/B sky130_fd_sc_hd__or2_4
X_19472_ _23324_/Q VGND VGND VPWR VPWR _19472_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16684_ _15918_/Y _23012_/A _15918_/Y _23012_/A VGND VGND VPWR VPWR _16688_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23937__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13896_ _13905_/A VGND VGND VPWR VPWR _13896_/X sky130_fd_sc_hd__buf_2
XFILLER_94_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18423_ _23813_/Q VGND VGND VPWR VPWR _18424_/D sky130_fd_sc_hd__inv_2
X_15635_ _15431_/X VGND VGND VPWR VPWR _15635_/X sky130_fd_sc_hd__buf_2
X_12847_ _25009_/Q VGND VGND VPWR VPWR _12878_/A sky130_fd_sc_hd__inv_2
XFILLER_64_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19156__B1 _19109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18354_ _24211_/Q _18491_/A _24217_/Q _18413_/A VGND VGND VPWR VPWR _18357_/C sky130_fd_sc_hd__a2bb2o_4
X_15566_ _15561_/X VGND VGND VPWR VPWR _15566_/X sky130_fd_sc_hd__buf_2
XANTENNA__16260__A1_N _14958_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12778_ _21980_/A VGND VGND VPWR VPWR _12778_/Y sky130_fd_sc_hd__inv_2
XPHY_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22745__A _24116_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _24004_/Q VGND VGND VPWR VPWR _17305_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14517_ _21752_/A _14517_/B VGND VGND VPWR VPWR _14517_/X sky130_fd_sc_hd__or2_4
X_11729_ _11728_/X VGND VGND VPWR VPWR _11729_/X sky130_fd_sc_hd__buf_2
X_18285_ _18273_/B VGND VGND VPWR VPWR _18286_/B sky130_fd_sc_hd__inv_2
X_15497_ HWDATA[15] VGND VGND VPWR VPWR _15497_/X sky130_fd_sc_hd__buf_2
XPHY_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17236_ _11596_/Y _17319_/A _11596_/Y _17319_/A VGND VGND VPWR VPWR _17236_/X sky130_fd_sc_hd__a2bb2o_4
X_14448_ _19904_/D _14448_/B VGND VGND VPWR VPWR _14448_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17558__B _17558_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15359__A _15358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11887__A _22006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17167_ _17086_/X _17161_/B _17166_/Y VGND VGND VPWR VPWR _24028_/D sky130_fd_sc_hd__and3_4
XANTENNA__24796__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14379_ _13429_/Y _14378_/Y VGND VGND VPWR VPWR _14380_/B sky130_fd_sc_hd__or2_4
XANTENNA__14940__B2 _24267_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16118_ _16116_/Y _16112_/X _15992_/X _16117_/X VGND VGND VPWR VPWR _24328_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16142__B1 _16141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24725__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17098_ _17097_/X VGND VGND VPWR VPWR _17099_/B sky130_fd_sc_hd__inv_2
XFILLER_116_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_151_0_HCLK clkbuf_7_75_0_HCLK/X VGND VGND VPWR VPWR _24372_/CLK sky130_fd_sc_hd__clkbuf_1
X_16049_ _16048_/Y _16046_/X _11522_/X _16046_/X VGND VGND VPWR VPWR _16049_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21096__A _21275_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19808_ _11635_/A VGND VGND VPWR VPWR _19808_/X sky130_fd_sc_hd__buf_2
XANTENNA__12511__A _12345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19739_ _22100_/B _19738_/X _19711_/X _19738_/X VGND VGND VPWR VPWR _23230_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15822__A _15414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22750_ _24347_/Q _22549_/A _22581_/X VGND VGND VPWR VPWR _22750_/X sky130_fd_sc_hd__o21a_4
XFILLER_53_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23678__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21701_ _22047_/A _19263_/A _19265_/A _21701_/D VGND VGND VPWR VPWR _21701_/X sky130_fd_sc_hd__or4_4
XANTENNA__21741__A2 _21300_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15956__B1 _15775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22681_ _22681_/A _22681_/B _22681_/C VGND VGND VPWR VPWR _22686_/B sky130_fd_sc_hd__and3_4
XANTENNA__21262__C _21193_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21742__A2_N _21408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24420_ _24590_/CLK _24420_/D HRESETn VGND VGND VPWR VPWR _24420_/Q sky130_fd_sc_hd__dfrtp_4
X_21632_ _21617_/A _21632_/B VGND VGND VPWR VPWR _21632_/X sky130_fd_sc_hd__or2_4
XFILLER_40_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24351_ _24333_/CLK _24351_/D HRESETn VGND VGND VPWR VPWR _16056_/A sky130_fd_sc_hd__dfrtp_4
X_21563_ _16544_/Y _21561_/X _15395_/Y _21562_/X VGND VGND VPWR VPWR _21564_/B sky130_fd_sc_hd__o22a_4
XANTENNA__15708__B1 _15286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17749__A _14577_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23302_ _23100_/CLK _19535_/X VGND VGND VPWR VPWR _19529_/A sky130_fd_sc_hd__dfxtp_4
X_20514_ _20512_/Y _20508_/X _20513_/X VGND VGND VPWR VPWR _20514_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15184__A1 _14941_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24282_ _24662_/CLK _24282_/D HRESETn VGND VGND VPWR VPWR _14901_/A sky130_fd_sc_hd__dfrtp_4
X_21494_ _15428_/X _21493_/X _23913_/Q _12063_/X VGND VGND VPWR VPWR _21494_/X sky130_fd_sc_hd__o22a_4
XFILLER_14_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23233_ _23401_/CLK _19729_/X VGND VGND VPWR VPWR _19726_/A sky130_fd_sc_hd__dfxtp_4
X_20445_ _20445_/A VGND VGND VPWR VPWR _20445_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22454__B1 _20750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24466__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23164_ _23332_/CLK _23164_/D VGND VGND VPWR VPWR _19910_/A sky130_fd_sc_hd__dfxtp_4
X_20376_ _20375_/X VGND VGND VPWR VPWR _20376_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12405__B _12534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22115_ _22083_/X _22114_/X _21062_/X VGND VGND VPWR VPWR _22138_/C sky130_fd_sc_hd__a21oi_4
XFILLER_133_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22206__B1 _14744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16684__B2 _23012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23095_ _23249_/CLK _23095_/D VGND VGND VPWR VPWR _23095_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_115_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22046_ _22046_/A _22042_/B VGND VGND VPWR VPWR _22046_/X sky130_fd_sc_hd__or2_4
XFILLER_0_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12421__A _12305_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22509__A1 _22879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23997_ _25214_/CLK _17384_/X HRESETn VGND VGND VPWR VPWR _17251_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13750_ _13769_/A _13769_/B _13716_/C _13716_/D VGND VGND VPWR VPWR _13757_/B sky130_fd_sc_hd__a211o_4
X_22948_ _14814_/Y _21544_/X _14920_/Y _22312_/B VGND VGND VPWR VPWR _22948_/X sky130_fd_sc_hd__o22a_4
X_12701_ _12701_/A _12701_/B VGND VGND VPWR VPWR _12704_/B sky130_fd_sc_hd__or2_4
XFILLER_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13681_ _13677_/C VGND VGND VPWR VPWR _13681_/X sky130_fd_sc_hd__buf_2
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_14_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_14_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_22879_ _22879_/A _22876_/X _22879_/C VGND VGND VPWR VPWR _22906_/A sky130_fd_sc_hd__and3_4
X_15420_ _22314_/B VGND VGND VPWR VPWR _16228_/A sky130_fd_sc_hd__buf_2
XFILLER_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12632_ _12632_/A _12632_/B _12632_/C _12631_/X VGND VGND VPWR VPWR _12632_/X sky130_fd_sc_hd__or4_4
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24618_ _24618_/CLK _15311_/X HRESETn VGND VGND VPWR VPWR _24618_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ _12651_/D _20822_/A _12651_/D _20822_/A VGND VGND VPWR VPWR _12563_/X sky130_fd_sc_hd__a2bb2o_4
X_15351_ _22696_/A _15345_/X _15350_/X _15345_/X VGND VGND VPWR VPWR _24605_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24549_ _24545_/CLK _24549_/D HRESETn VGND VGND VPWR VPWR _24549_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16563__A _20863_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11514_ _11514_/A _14020_/A VGND VGND VPWR VPWR _11514_/X sky130_fd_sc_hd__or2_4
X_14302_ _24785_/Q VGND VGND VPWR VPWR _14302_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11984__B2 _11965_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18070_ _18068_/X _11746_/Y _18069_/X VGND VGND VPWR VPWR _19467_/A sky130_fd_sc_hd__or3_4
XFILLER_106_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ _12418_/C _12409_/X VGND VGND VPWR VPWR _12495_/B sky130_fd_sc_hd__or2_4
X_15282_ _15282_/A VGND VGND VPWR VPWR _15282_/X sky130_fd_sc_hd__buf_2
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17021_ _17021_/A VGND VGND VPWR VPWR _17021_/Y sky130_fd_sc_hd__inv_2
X_14233_ _14230_/Y _14226_/X _14232_/X _14226_/X VGND VGND VPWR VPWR _14233_/X sky130_fd_sc_hd__a2bb2o_4
X_14164_ _14168_/A VGND VGND VPWR VPWR _14165_/B sky130_fd_sc_hd__buf_2
XFILLER_67_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16124__B1 _15709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20235__D _20235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20813__A _15455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15478__A2 _15461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13115_ _11711_/X _13088_/X _13113_/X _25003_/Q _13114_/X VGND VGND VPWR VPWR _13115_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__24136__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_224_0_HCLK clkbuf_8_225_0_HCLK/A VGND VGND VPWR VPWR _24042_/CLK sky130_fd_sc_hd__clkbuf_1
X_14095_ _14093_/Y _14091_/X _14094_/X _14091_/X VGND VGND VPWR VPWR _14095_/X sky130_fd_sc_hd__a2bb2o_4
X_18972_ _13068_/B VGND VGND VPWR VPWR _18972_/Y sky130_fd_sc_hd__inv_2
X_13046_ _13049_/A _23598_/Q VGND VGND VPWR VPWR _13047_/C sky130_fd_sc_hd__or2_4
X_17923_ _17955_/A _17923_/B _17923_/C VGND VGND VPWR VPWR _17923_/X sky130_fd_sc_hd__and3_4
XFILLER_79_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17854_ _17780_/A _17852_/X _17853_/X VGND VGND VPWR VPWR _17858_/B sky130_fd_sc_hd__and3_4
XFILLER_61_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16805_ _15902_/Y _24062_/Q _24396_/Q _16921_/C VGND VGND VPWR VPWR _16809_/A sky130_fd_sc_hd__a2bb2o_4
X_17785_ _17739_/A _17785_/B _17785_/C VGND VGND VPWR VPWR _17785_/X sky130_fd_sc_hd__and3_4
X_14997_ _14997_/A _14997_/B VGND VGND VPWR VPWR _14997_/X sky130_fd_sc_hd__or2_4
XFILLER_81_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19524_ _19522_/Y _19523_/X _19459_/X _19523_/X VGND VGND VPWR VPWR _19524_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15642__A _15637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16736_ _15935_/Y _22853_/A _24380_/Q _17497_/D VGND VGND VPWR VPWR _16739_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21363__B _11986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13948_ _14247_/A _13937_/X _13938_/X _13947_/Y VGND VGND VPWR VPWR _24895_/D sky130_fd_sc_hd__o22a_4
XFILLER_75_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23771__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_1_1_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19455_ _19455_/A VGND VGND VPWR VPWR _19455_/X sky130_fd_sc_hd__buf_2
X_16667_ _14699_/Y _16663_/X _16373_/X _16666_/X VGND VGND VPWR VPWR _16667_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23700__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13879_ _13842_/X _13879_/B VGND VGND VPWR VPWR _13887_/A sky130_fd_sc_hd__or2_4
X_18406_ _18402_/X _18403_/X _18404_/X _18405_/X VGND VGND VPWR VPWR _18406_/X sky130_fd_sc_hd__or4_4
X_15618_ _15611_/X _15617_/X _15505_/X _24514_/Q _15612_/X VGND VGND VPWR VPWR _24514_/D
+ sky130_fd_sc_hd__a32o_4
X_19386_ _19372_/Y VGND VGND VPWR VPWR _19386_/X sky130_fd_sc_hd__buf_2
X_16598_ _16581_/X _16597_/X _11585_/A _24139_/Q _16590_/X VGND VGND VPWR VPWR _16598_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18337_ _18336_/X VGND VGND VPWR VPWR _23845_/D sky130_fd_sc_hd__inv_2
XFILLER_37_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15549_ _19452_/A VGND VGND VPWR VPWR _15549_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22684__B1 _20777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24977__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18268_ _18268_/A _18268_/B VGND VGND VPWR VPWR _18269_/C sky130_fd_sc_hd__or2_4
XANTENNA__24906__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15705__A3 _15704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17219_ _20735_/A VGND VGND VPWR VPWR _17219_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18199_ _18199_/A VGND VGND VPWR VPWR _18242_/A sky130_fd_sc_hd__inv_2
Xclkbuf_6_34_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_34_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20230_ _20225_/X _20229_/X VGND VGND VPWR VPWR _20230_/X sky130_fd_sc_hd__or2_4
XFILLER_128_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16115__B1 _15897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21819__A _20979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15469__A2 _15461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20161_ _20192_/A _20160_/Y VGND VGND VPWR VPWR _20161_/X sky130_fd_sc_hd__and2_4
XANTENNA__21538__B _21458_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22739__A1 _16501_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22739__B2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20092_ _21142_/B _20089_/X _19617_/A _20089_/X VGND VGND VPWR VPWR _23095_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13337__A _13337_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23920_ _24757_/CLK _23920_/D HRESETn VGND VGND VPWR VPWR _23920_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23859__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19537__A2_N _19534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21554__A _21860_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23851_ _23845_/CLK _18320_/X HRESETn VGND VGND VPWR VPWR _23851_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22802_ _24118_/Q _22745_/B VGND VGND VPWR VPWR _22805_/B sky130_fd_sc_hd__or2_4
X_20994_ _20994_/A VGND VGND VPWR VPWR _21006_/A sky130_fd_sc_hd__buf_2
X_23782_ _24980_/CLK _13494_/Y HRESETn VGND VGND VPWR VPWR _14106_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__22911__A1 _21490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22911__B2 _22840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22733_ _24417_/Q _22281_/X _20782_/A _22732_/X VGND VGND VPWR VPWR _22734_/C sky130_fd_sc_hd__a211o_4
XFILLER_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13072__A _13065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22664_ _21540_/X _22662_/X _20839_/X _22663_/X VGND VGND VPWR VPWR _22664_/X sky130_fd_sc_hd__o22a_4
XFILLER_129_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22385__A _22385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21615_ _21612_/A _21615_/B VGND VGND VPWR VPWR _21615_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_116_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_233_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24403_ _24620_/CLK _15888_/X HRESETn VGND VGND VPWR VPWR _24403_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17479__A _16710_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22595_ _22595_/A _21979_/X VGND VGND VPWR VPWR _22595_/X sky130_fd_sc_hd__or2_4
XFILLER_103_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21546_ _15578_/B VGND VGND VPWR VPWR _21546_/X sky130_fd_sc_hd__buf_2
XANTENNA__24647__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24334_ _24222_/CLK _16103_/X HRESETn VGND VGND VPWR VPWR _16102_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19694__A _19688_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24265_ _24264_/CLK _16280_/X HRESETn VGND VGND VPWR VPWR _14897_/A sky130_fd_sc_hd__dfrtp_4
X_21477_ _21340_/A _21477_/B VGND VGND VPWR VPWR _21477_/X sky130_fd_sc_hd__or2_4
XANTENNA__12416__A _12416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22832__B _22813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23216_ _23401_/CLK _23216_/D VGND VGND VPWR VPWR _19774_/A sky130_fd_sc_hd__dfxtp_4
X_20428_ _20428_/A VGND VGND VPWR VPWR _20428_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16106__B1 _15978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24196_ _24192_/CLK _16461_/X HRESETn VGND VGND VPWR VPWR _24196_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23147_ _23596_/CLK _19956_/X VGND VGND VPWR VPWR _19955_/A sky130_fd_sc_hd__dfxtp_4
X_20359_ _17174_/A _17174_/B VGND VGND VPWR VPWR _20359_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__21448__B _21448_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23078_ _23109_/CLK _23078_/D VGND VGND VPWR VPWR _23078_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13340__B1 _11612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14920_ _24284_/Q VGND VGND VPWR VPWR _14920_/Y sky130_fd_sc_hd__inv_2
X_22029_ _21544_/A VGND VGND VPWR VPWR _22029_/X sky130_fd_sc_hd__buf_2
XFILLER_121_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17942__A _14577_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_54_0_HCLK clkbuf_8_55_0_HCLK/A VGND VGND VPWR VPWR _23957_/CLK sky130_fd_sc_hd__clkbuf_1
X_14851_ _24706_/Q _14850_/Y _24706_/Q _14850_/Y VGND VGND VPWR VPWR _14855_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16558__A _13644_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13802_ _13866_/A VGND VGND VPWR VPWR _13833_/A sky130_fd_sc_hd__buf_2
XFILLER_112_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15632__A2 _15617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15462__A _13357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17570_ _17497_/B _17548_/X VGND VGND VPWR VPWR _17570_/X sky130_fd_sc_hd__or2_4
X_14782_ _24702_/Q VGND VGND VPWR VPWR _15022_/A sky130_fd_sc_hd__inv_2
X_11994_ _25145_/Q VGND VGND VPWR VPWR _11994_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22902__A1 _16693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16521_ _16520_/Y _16518_/X _15369_/X _16518_/X VGND VGND VPWR VPWR _16521_/X sky130_fd_sc_hd__a2bb2o_4
X_13733_ _13730_/A _24637_/Q _13726_/X _13732_/B VGND VGND VPWR VPWR _13734_/A sky130_fd_sc_hd__or4_4
XANTENNA__19869__A _19876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14078__A _16559_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19240_ _19234_/Y _19239_/X _11835_/X _19239_/X VGND VGND VPWR VPWR _23406_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16452_ _16452_/A VGND VGND VPWR VPWR _16452_/X sky130_fd_sc_hd__buf_2
XFILLER_31_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13664_ _13434_/Y _13661_/X _13663_/X _13661_/X VGND VGND VPWR VPWR _13664_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16593__B1 _16179_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20808__A _20808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15403_ _24585_/Q VGND VGND VPWR VPWR _15403_/Y sky130_fd_sc_hd__inv_2
X_12615_ _24530_/Q VGND VGND VPWR VPWR _12615_/Y sky130_fd_sc_hd__inv_2
X_19171_ _19166_/Y _19169_/X _19170_/X _19169_/X VGND VGND VPWR VPWR _19171_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17389__A _17270_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16383_ _16383_/A VGND VGND VPWR VPWR _16383_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22666__B1 _17497_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ _13559_/X _13593_/Y _13594_/X _13587_/X _11657_/A VGND VGND VPWR VPWR _24953_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18122_ _23881_/Q VGND VGND VPWR VPWR _18122_/Y sky130_fd_sc_hd__inv_2
X_15334_ _15331_/Y _15327_/X _15332_/X _15333_/X VGND VGND VPWR VPWR _15334_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24388__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12546_ _24508_/Q VGND VGND VPWR VPWR _12546_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18053_ _20034_/A _18052_/X _20034_/A _18052_/X VGND VGND VPWR VPWR _18053_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24317__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15265_ _13722_/X _15260_/X _15256_/X _24637_/Q _15262_/X VGND VGND VPWR VPWR _15265_/X
+ sky130_fd_sc_hd__a32o_4
X_12477_ _12474_/C _12466_/B VGND VGND VPWR VPWR _12478_/B sky130_fd_sc_hd__or2_4
X_17004_ _17000_/X _17001_/X _17004_/C _17003_/X VGND VGND VPWR VPWR _17004_/X sky130_fd_sc_hd__or4_4
X_14216_ _14215_/Y _14212_/X _14094_/X _14201_/X VGND VGND VPWR VPWR _24818_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_6_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15196_ _15224_/A _15110_/B _15112_/C _15229_/A VGND VGND VPWR VPWR _15197_/B sky130_fd_sc_hd__or4_4
XFILLER_125_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14147_ _14147_/A VGND VGND VPWR VPWR _14147_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14078_ _16559_/A _17197_/B VGND VGND VPWR VPWR _14079_/A sky130_fd_sc_hd__nor2_4
X_18955_ _17871_/B VGND VGND VPWR VPWR _18955_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13331__B1 _13330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13029_ _13042_/A VGND VGND VPWR VPWR _13049_/A sky130_fd_sc_hd__buf_2
X_17906_ _16022_/Y _17898_/X _17905_/X VGND VGND VPWR VPWR _17906_/X sky130_fd_sc_hd__and3_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18886_ _23531_/Q VGND VGND VPWR VPWR _18886_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23952__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21374__A _21374_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25176__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17837_ _17742_/A VGND VGND VPWR VPWR _17934_/A sky130_fd_sc_hd__buf_2
XFILLER_120_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25105__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21093__B _21093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17768_ _17708_/X _17766_/X _23932_/Q _17767_/X VGND VGND VPWR VPWR _17768_/X sky130_fd_sc_hd__o22a_4
XFILLER_130_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16719_ _15957_/A _17558_/B _15989_/Y _23947_/Q VGND VGND VPWR VPWR _16719_/X sky130_fd_sc_hd__a2bb2o_4
X_19507_ _19505_/Y _19501_/X _19506_/X _19488_/Y VGND VGND VPWR VPWR _23311_/D sky130_fd_sc_hd__a2bb2o_4
X_17699_ _17676_/X _17697_/X _17699_/C VGND VGND VPWR VPWR _17699_/X sky130_fd_sc_hd__and3_4
X_19438_ _23334_/Q VGND VGND VPWR VPWR _19438_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19369_ _19368_/Y _19363_/X _19232_/X _19349_/Y VGND VGND VPWR VPWR _23359_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21400_ _21400_/A VGND VGND VPWR VPWR _21400_/X sky130_fd_sc_hd__buf_2
X_22380_ _22360_/X _22363_/X _22368_/X _22375_/X _22379_/X VGND VGND VPWR VPWR _22380_/X
+ sky130_fd_sc_hd__o41a_4
XANTENNA__12070__B1 _11643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20132__A1 _23077_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24740__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19010__C _14482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21331_ _21327_/X _21330_/X _18049_/X VGND VGND VPWR VPWR _21331_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24058__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21880__A1 _15271_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24050_ _24049_/CLK _17090_/X HRESETn VGND VGND VPWR VPWR _17089_/A sky130_fd_sc_hd__dfrtp_4
X_21262_ _21262_/A _21128_/X _21193_/X _21261_/X VGND VGND VPWR VPWR HRDATA[1] sky130_fd_sc_hd__or4_4
XFILLER_89_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23001_ _22968_/A _23001_/B VGND VGND VPWR VPWR _23001_/X sky130_fd_sc_hd__and2_4
X_20213_ _14102_/X VGND VGND VPWR VPWR _20225_/B sky130_fd_sc_hd__inv_2
X_21193_ _21176_/Y _21190_/Y _21192_/X VGND VGND VPWR VPWR _21193_/X sky130_fd_sc_hd__o21a_4
XFILLER_104_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20144_ _20143_/Y _20141_/X _15520_/X _20141_/X VGND VGND VPWR VPWR _20144_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17762__A _14569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20075_ _19530_/X _19282_/B _19531_/X VGND VGND VPWR VPWR _20076_/A sky130_fd_sc_hd__or3_4
X_24952_ _24757_/CLK _13597_/X HRESETn VGND VGND VPWR VPWR _11670_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23693__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23903_ _23356_/CLK _18032_/X HRESETn VGND VGND VPWR VPWR _23903_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23622__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24883_ _24884_/CLK _24883_/D HRESETn VGND VGND VPWR VPWR _13925_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_57_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23834_ _23830_/CLK _18492_/X HRESETn VGND VGND VPWR VPWR _23834_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21148__B1 _17639_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19689__A _19688_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20977_ _20971_/A VGND VGND VPWR VPWR _20978_/A sky130_fd_sc_hd__buf_2
XFILLER_72_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24899__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23765_ _23767_/CLK _20266_/X HRESETn VGND VGND VPWR VPWR _23765_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17367__A2 _17366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24828__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22716_ _22712_/X _22716_/B _22716_/C _22715_/X VGND VGND VPWR VPWR _22716_/X sky130_fd_sc_hd__or4_4
X_23696_ _24161_/CLK _20424_/Y HRESETn VGND VGND VPWR VPWR _13499_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22648__B1 _24414_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22647_ _22992_/B VGND VGND VPWR VPWR _22647_/X sky130_fd_sc_hd__buf_2
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12400_ _25098_/Q VGND VGND VPWR VPWR _12401_/B sky130_fd_sc_hd__inv_2
X_13380_ _13391_/A _13377_/X _11981_/X _13377_/X VGND VGND VPWR VPWR _13380_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24481__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16327__B1 _16251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22578_ _24143_/Q _15692_/A _22576_/X _22577_/X VGND VGND VPWR VPWR _22579_/C sky130_fd_sc_hd__a211o_4
XFILLER_127_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12331_ _25094_/Q VGND VGND VPWR VPWR _12448_/A sky130_fd_sc_hd__inv_2
XANTENNA__24410__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24317_ _24319_/CLK _24317_/D HRESETn VGND VGND VPWR VPWR _24317_/Q sky130_fd_sc_hd__dfrtp_4
X_21529_ _21245_/X VGND VGND VPWR VPWR _21529_/X sky130_fd_sc_hd__buf_2
XANTENNA__12146__A _24565_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12262_ _12127_/Y _12257_/B _12259_/B _12195_/X VGND VGND VPWR VPWR _12262_/X sky130_fd_sc_hd__a211o_4
X_15050_ _15019_/B _15049_/X VGND VGND VPWR VPWR _15051_/A sky130_fd_sc_hd__or2_4
X_24248_ _24213_/CLK _16322_/X HRESETn VGND VGND VPWR VPWR _16320_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14001_ _13997_/Y _14000_/Y _13992_/X VGND VGND VPWR VPWR _14001_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15457__A _15414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12193_ _12193_/A _12193_/B VGND VGND VPWR VPWR _12193_/X sky130_fd_sc_hd__or2_4
X_24179_ _24112_/CLK _24179_/D HRESETn VGND VGND VPWR VPWR _24179_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14105__A2 _14100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17094__D _17124_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22179__A2 _21178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18740_ _18739_/X VGND VGND VPWR VPWR _18740_/X sky130_fd_sc_hd__buf_2
X_15952_ _22639_/A VGND VGND VPWR VPWR _15952_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14903_ _24650_/Q VGND VGND VPWR VPWR _14903_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18671_ _18670_/Y _18668_/X _17202_/X _18668_/X VGND VGND VPWR VPWR _23605_/D sky130_fd_sc_hd__a2bb2o_4
X_15883_ _15882_/Y _15880_/X _15788_/X _15880_/X VGND VGND VPWR VPWR _24405_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17622_ _20778_/A _17622_/B VGND VGND VPWR VPWR _17622_/X sky130_fd_sc_hd__or2_4
XFILLER_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12311__A1_N _12451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14834_ _15034_/A _24142_/Q _14712_/X _14833_/Y VGND VGND VPWR VPWR _14834_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16612__A1_N _14801_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14813__B1 _15033_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17553_ _16692_/A _17553_/B VGND VGND VPWR VPWR _17553_/X sky130_fd_sc_hd__or2_4
XANTENNA__11627__B1 _11626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21922__A _20968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14765_ _24705_/Q VGND VGND VPWR VPWR _14765_/Y sky130_fd_sc_hd__inv_2
X_11977_ _25150_/Q VGND VGND VPWR VPWR _11977_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16504_ _22695_/A _16499_/X _16334_/X _16499_/X VGND VGND VPWR VPWR _24179_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13716_ _13716_/A _13716_/B _13716_/C _13716_/D VGND VGND VPWR VPWR _13716_/X sky130_fd_sc_hd__or4_4
X_17484_ _23946_/Q VGND VGND VPWR VPWR _17484_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24569__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14696_ _15064_/A _16658_/A _15064_/A _16658_/A VGND VGND VPWR VPWR _14696_/X sky130_fd_sc_hd__a2bb2o_4
X_19223_ _19223_/A VGND VGND VPWR VPWR _19223_/Y sky130_fd_sc_hd__inv_2
X_16435_ _16432_/Y _16434_/X _16179_/X _16434_/X VGND VGND VPWR VPWR _24206_/D sky130_fd_sc_hd__a2bb2o_4
X_13647_ _12065_/A _13611_/X VGND VGND VPWR VPWR _13647_/Y sky130_fd_sc_hd__nor2_4
XFILLER_73_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19154_ _19151_/Y _19146_/X _19152_/X _19153_/X VGND VGND VPWR VPWR _19154_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16366_ _16366_/A VGND VGND VPWR VPWR _16366_/Y sky130_fd_sc_hd__inv_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ _11653_/A _13566_/B VGND VGND VPWR VPWR _13578_/X sky130_fd_sc_hd__or2_4
XANTENNA__14967__A2_N _24285_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18105_ _18097_/X _18104_/Y _18089_/A _18096_/Y VGND VGND VPWR VPWR _23888_/D sky130_fd_sc_hd__a2bb2o_4
X_15317_ _21019_/A VGND VGND VPWR VPWR _20926_/A sky130_fd_sc_hd__buf_2
XANTENNA__24151__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12529_ _12405_/D _12423_/A VGND VGND VPWR VPWR _12536_/B sky130_fd_sc_hd__or2_4
X_19085_ _19083_/Y _19079_/X _19041_/X _19084_/X VGND VGND VPWR VPWR _23460_/D sky130_fd_sc_hd__a2bb2o_4
X_16297_ _16296_/Y VGND VGND VPWR VPWR _18263_/A sky130_fd_sc_hd__buf_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18036_ _18023_/X _18033_/X _18035_/Y VGND VGND VPWR VPWR _18036_/X sky130_fd_sc_hd__o21a_4
X_15248_ _13761_/A _15247_/X _15240_/X _13776_/C _15245_/X VGND VGND VPWR VPWR _24647_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12355__B2 _24472_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22811__B1 _21562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15179_ _15179_/A _15183_/B VGND VGND VPWR VPWR _15180_/C sky130_fd_sc_hd__nand2_4
XFILLER_126_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19987_ _19986_/Y _19982_/X _19859_/A _19982_/A VGND VGND VPWR VPWR _19987_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18678__A HWDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18938_ _18801_/X VGND VGND VPWR VPWR _18938_/X sky130_fd_sc_hd__buf_2
XFILLER_100_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
.ends

