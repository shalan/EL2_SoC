
`default_nettype none
`timescale 1ns/1ns
//`define		USE_DFFRAM_BEH

module soc_core (
	input HCLK, 
	input HRESETn,
	
	input wire 			NMI,
	input wire [7:0]	SYSTICKCLKDIV,

	input wire  [3: 0] 	fdi_Sys0_S0,
	output wire [3: 0] 	fdo_Sys0_S0,
	output wire [0: 0] 	fdoe_Sys0_S0,
	output wire [0: 0] 	fsclk_Sys0_S0,
	output wire [0: 0] 	fcen_Sys0_S0,

	input wire  [15: 0] GPIOIN_Sys0_S2,
	output wire [15: 0] GPIOOUT_Sys0_S2,
	output wire [15: 0] GPIOPU_Sys0_S2,
	output wire [15: 0] GPIOPD_Sys0_S2,
	output wire [15: 0] GPIOOEN_Sys0_S2,

	input wire [0: 0] RsRx_Sys0_SS0_S0,
	output wire [0: 0] RsTx_Sys0_SS0_S0,

	input wire [0: 0] RsRx_Sys0_SS0_S1,
	output wire [0: 0] RsTx_Sys0_SS0_S1,

	input wire [0: 0] MSI_Sys0_SS0_S2,
	output wire [0: 0] MSO_Sys0_SS0_S2,
	output wire [0: 0] SSn_Sys0_SS0_S2,
	output wire [0: 0] SCLK_Sys0_SS0_S2,
	input wire [0: 0] MSI_Sys0_SS0_S3,
	output wire [0: 0] MSO_Sys0_SS0_S3,
	output wire [0: 0] SSn_Sys0_SS0_S3,
	output wire [0: 0] SCLK_Sys0_SS0_S3,
	input wire [0: 0] scl_i_Sys0_SS0_S4,
	output wire [0: 0] scl_o_Sys0_SS0_S4,
	output wire [0: 0] scl_oen_o_Sys0_SS0_S4,
	input wire [0: 0] sda_i_Sys0_SS0_S4,
	output wire [0: 0] sda_o_Sys0_SS0_S4,
	output wire [0: 0] sda_oen_o_Sys0_SS0_S4,

	input wire [0: 0] scl_i_Sys0_SS0_S5,
	output wire [0: 0] scl_o_Sys0_SS0_S5,
	output wire [0: 0] scl_oen_o_Sys0_SS0_S5,
	input wire [0: 0] sda_i_Sys0_SS0_S5,
	output wire [0: 0] sda_o_Sys0_SS0_S5,
	output wire [0: 0] sda_oen_o_Sys0_SS0_S5,

	output wire [0: 0] pwm_Sys0_SS0_S6,
	output wire [0: 0] pwm_Sys0_SS0_S7
);

	wire [`AW-1: 0] HADDR_Sys0;
	wire [`DW-1: 0] HWDATA_Sys0;
	wire HWRITE_Sys0;
	wire [1: 0] HTRANS_Sys0;
	wire [2:0] HSIZE_Sys0;

	wire HREADY_Sys0;
	wire [`DW-1: 0] HRDATA_Sys0;

	wire [`DW-1: 0] SRAMRDATA_Sys0_S1;
	wire [7: 0] SRAMWEN_Sys0_S1;
	wire [`DW-1: 0] SRAMWDATA_Sys0_S1;
	wire [0: 0] SRAMCS0_Sys0_S1;
	wire [9: 0] SRAMADDR_Sys0_S1;

	// AHB LITE Master2 Signals
	wire [`AW-1:0] M0_HADDR, M1_HADDR;
	wire [0:0] M0_HREADY, M1_HREADY;
	wire [0:0] M0_HWRITE, M1_HWRITE;
	wire [1:0] M0_HTRANS, M1_HTRANS;
	wire [2:0] M0_HSIZE, M1_HSIZE;
	wire [`DW-1:0] M0_HWDATA, M1_HWDATA;
	wire [`DW-1:0] M0_HRDATA, M1_HRDATA;
	
	wire [31: 0] M0_IRQ;

	wire [3:0] M0_HPROT, M1_HPROT;
	wire [2:0] M0_HBURST, M1_HBURST;
	wire M0_HMASTLOCK,  M1_HMASTLOCK;

	wire M0_HBUSREQ, M1_HBUSREQ;
	wire M0_HLOCK;
	wire M0_HGRANT, M1_HGRANT;

	assign M0_HRDATA = HRDATA_Sys0;
	assign M1_HRDATA = HRDATA_Sys0;

	assign HADDR_Sys0 = M0_HADDR; 
	assign HWDATA_Sys0 = M0_HWDATA; 
	assign HWRITE_Sys0 = M0_HWRITE; 
	assign HTRANS_Sys0 = M0_HTRANS; 
	assign HSIZE_Sys0 = M0_HSIZE;

	//AHBlite_SYS0 instantiation
	AHBlite_sys_0 ahb_sys_0_uut(

		.HCLK(HCLK),
		.HRESETn(HRESETn),
         
		.M0_HADDR(HADDR_Sys0),
		.M0_HWDATA(HWDATA_Sys0),
		.M0_HWRITE(HWRITE_Sys0),
		.M0_HTRANS(HTRANS_Sys0),
		.M0_HSIZE(HSIZE_Sys0),
		.M0_HBURST(M0_HBURST),
		.M0_HPROT(M0_HPROT),
		.M0_HMASTLOCK(M0_HMASTLOCK),
		.M0_HBUSREQ(M0_HBUSREQ),
		.M0_HGRANT(M0_HGRANT),
		.M0_HREADY(M0_HREADY),

		.M1_HADDR(M1_HADDR),
		.M1_HWDATA(M1_HWDATA),
		.M1_HWRITE(M1_HWRITE),
		.M1_HTRANS(M1_HTRANS),
		.M1_HSIZE(M1_HSIZE),
		.M1_HBURST(M1_HBURST),
		.M1_HPROT(M1_HPROT),
		.M1_HMASTLOCK(M1_HMASTLOCK),
		.M1_HBUSREQ(M1_HBUSREQ),
		.M1_HGRANT(M1_HGRANT),
		.M1_HREADY(M1_HREADY),

		.HRDATA(HRDATA_Sys0),
		
		// QSPI Interface
		.fdi_S0(fdi_Sys0_S0),
		.fdo_S0(fdo_Sys0_S0),
		.fdoe_S0(fdoe_Sys0_S0),
		.fsclk_S0(fsclk_Sys0_S0),
		.fcen_S0(fcen_Sys0_S0),

		// SRAM Interface
		.SRAMRDATA_S1(SRAMRDATA_Sys0_S1),
		.SRAMWEN_S1(SRAMWEN_Sys0_S1),
		.SRAMWDATA_S1(SRAMWDATA_Sys0_S1),
		.SRAMCS0_S1(SRAMCS0_Sys0_S1),
		.SRAMADDR_S1(SRAMADDR_Sys0_S1),

		// GPIO Interface
		.GPIOIN_S2(GPIOIN_Sys0_S2),
		.GPIOOUT_S2(GPIOOUT_Sys0_S2),
		.GPIOPU_S2(GPIOPU_Sys0_S2),
		.GPIOPD_S2(GPIOPD_Sys0_S2),
		.GPIOOEN_S2(GPIOOEN_Sys0_S2),
		
		// APB Bus
		// UART 0
		.RsRx_SS0_S0(RsRx_Sys0_SS0_S0),
		.RsTx_SS0_S0(RsTx_Sys0_SS0_S0),
		
		// UART 1
		.RsRx_SS0_S1(RsRx_Sys0_SS0_S1),
		.RsTx_SS0_S1(RsTx_Sys0_SS0_S1),

		// SPI 0 Interface
		.MSI_SS0_S2(MSI_Sys0_SS0_S2),
		.MSO_SS0_S2(MSO_Sys0_SS0_S2),
		.SSn_SS0_S2(SSn_Sys0_SS0_S2),
		.SCLK_SS0_S2(SCLK_Sys0_SS0_S2),

		// SPI 1 Interface
		.MSI_SS0_S3(MSI_Sys0_SS0_S3),
		.MSO_SS0_S3(MSO_Sys0_SS0_S3),
		.SSn_SS0_S3(SSn_Sys0_SS0_S3),
		.SCLK_SS0_S3(SCLK_Sys0_SS0_S3),

		// I2C 0 Interface
		.scl_i_SS0_S4(scl_i_Sys0_SS0_S4),
		.scl_o_SS0_S4(scl_o_Sys0_SS0_S4),
		.scl_oen_o_SS0_S4(scl_oen_o_Sys0_SS0_S4),
		.sda_i_SS0_S4(sda_i_Sys0_SS0_S4),
		.sda_o_SS0_S4(sda_o_Sys0_SS0_S4),
		.sda_oen_o_SS0_S4(sda_oen_o_Sys0_SS0_S4),

		// I2C 1 Interface
		.scl_i_SS0_S5(scl_i_Sys0_SS0_S5),
		.scl_o_SS0_S5(scl_o_Sys0_SS0_S5),
		.scl_oen_o_SS0_S5(scl_oen_o_Sys0_SS0_S5),
		.sda_i_SS0_S5(sda_i_Sys0_SS0_S5),
		.sda_o_SS0_S5(sda_o_Sys0_SS0_S5),
		.sda_oen_o_SS0_S5(sda_oen_o_Sys0_SS0_S5),

		// PMW 0 & 1 Interfaces
		.pwm_SS0_S6(pwm_Sys0_SS0_S6),
		.pwm_SS0_S7(pwm_Sys0_SS0_S7),

		.IRQ(M0_IRQ)

	);


	RAM_1024x64 RAM (
		.CLK(HCLK),
		.WE(SRAMWEN_Sys0_S1),
		.EN(SRAMCS0_Sys0_S1),
		.Di(SRAMWDATA_Sys0_S1),
		.Do(SRAMRDATA_Sys0_S1),
		.A(SRAMADDR_Sys0_S1[9:0])
	);

	// Instantiation of NfiVe32
	el2_n5_soc_wrapper EL2 (
		.HCLK(HCLK),
		.HRESETn(HRESETn),
		
		// Instructions
		.M0_HADDR(M0_HADDR),
		.M0_HREADY(M0_HREADY),
		.M0_HWRITE(M0_HWRITE),
		.M0_HTRANS(M0_HTRANS),
		.M0_HSIZE(M0_HSIZE),
		.M0_HWDATA(M0_HWDATA),
		.M0_HRDATA(M0_HRDATA),
		.M0_HBURST(M0_HBURST),
		.M0_HPROT(M0_HPROT),
		.M0_HMASTLOCK(M0_HMASTLOCK),
		.M0_HGRANT(M0_HGRANT),
		.M0_HBUSREQ(M0_HBUSREQ),

		// LSU
		.M1_HADDR(M1_HADDR),
		.M1_HREADY(M1_HREADY),
		.M1_HWRITE(M1_HWRITE),
		.M1_HTRANS(M1_HTRANS),
		.M1_HSIZE(M1_HSIZE),
		.M1_HWDATA(M1_HWDATA),
		.M1_HRDATA(M1_HRDATA),
		.M1_HBURST(M1_HBURST),
		.M1_HPROT(M1_HPROT),
		.M1_HMASTLOCK(M1_HMASTLOCK),
		.M1_HGRANT(M1_HGRANT),
		.M1_HBUSREQ(M1_HBUSREQ),

		//NMI
		.NMI(NMI),

		//Interrupts
		.IRQ(M0_IRQ[14:0]),

		// SYSTICK Divisor
		.SYSTICKCLKDIV(SYSTICKCLKDIV)
	);
  endmodule
  