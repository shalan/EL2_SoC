magic
tech sky130A
magscale 1 2
timestamp 1611408210
<< obsli1 >>
rect 949 2159 278852 297585
<< obsm1 >>
rect 14 8 279390 298172
<< metal2 >>
rect 478 0 534 800
rect 1490 0 1546 800
rect 2594 0 2650 800
rect 3698 0 3754 800
rect 4710 0 4766 800
rect 5814 0 5870 800
rect 6918 0 6974 800
rect 8022 0 8078 800
rect 9034 0 9090 800
rect 10138 0 10194 800
rect 11242 0 11298 800
rect 12346 0 12402 800
rect 13358 0 13414 800
rect 14462 0 14518 800
rect 15566 0 15622 800
rect 16670 0 16726 800
rect 17682 0 17738 800
rect 18786 0 18842 800
rect 19890 0 19946 800
rect 20994 0 21050 800
rect 22006 0 22062 800
rect 23110 0 23166 800
rect 24214 0 24270 800
rect 25318 0 25374 800
rect 26330 0 26386 800
rect 27434 0 27490 800
rect 28538 0 28594 800
rect 29642 0 29698 800
rect 30654 0 30710 800
rect 31758 0 31814 800
rect 32862 0 32918 800
rect 33966 0 34022 800
rect 34978 0 35034 800
rect 36082 0 36138 800
rect 37186 0 37242 800
rect 38290 0 38346 800
rect 39302 0 39358 800
rect 40406 0 40462 800
rect 41510 0 41566 800
rect 42614 0 42670 800
rect 43626 0 43682 800
rect 44730 0 44786 800
rect 45834 0 45890 800
rect 46938 0 46994 800
rect 47950 0 48006 800
rect 49054 0 49110 800
rect 50158 0 50214 800
rect 51262 0 51318 800
rect 52274 0 52330 800
rect 53378 0 53434 800
rect 54482 0 54538 800
rect 55586 0 55642 800
rect 56598 0 56654 800
rect 57702 0 57758 800
rect 58806 0 58862 800
rect 59910 0 59966 800
rect 60922 0 60978 800
rect 62026 0 62082 800
rect 63130 0 63186 800
rect 64234 0 64290 800
rect 65246 0 65302 800
rect 66350 0 66406 800
rect 67454 0 67510 800
rect 68558 0 68614 800
rect 69570 0 69626 800
rect 70674 0 70730 800
rect 71778 0 71834 800
rect 72882 0 72938 800
rect 73894 0 73950 800
rect 74998 0 75054 800
rect 76102 0 76158 800
rect 77206 0 77262 800
rect 78218 0 78274 800
rect 79322 0 79378 800
rect 80426 0 80482 800
rect 81530 0 81586 800
rect 82542 0 82598 800
rect 83646 0 83702 800
rect 84750 0 84806 800
rect 85854 0 85910 800
rect 86866 0 86922 800
rect 87970 0 88026 800
rect 89074 0 89130 800
rect 90178 0 90234 800
rect 91190 0 91246 800
rect 92294 0 92350 800
rect 93398 0 93454 800
rect 94502 0 94558 800
rect 95514 0 95570 800
rect 96618 0 96674 800
rect 97722 0 97778 800
rect 98826 0 98882 800
rect 99838 0 99894 800
rect 100942 0 100998 800
rect 102046 0 102102 800
rect 103150 0 103206 800
rect 104162 0 104218 800
rect 105266 0 105322 800
rect 106370 0 106426 800
rect 107474 0 107530 800
rect 108486 0 108542 800
rect 109590 0 109646 800
rect 110694 0 110750 800
rect 111798 0 111854 800
rect 112810 0 112866 800
rect 113914 0 113970 800
rect 115018 0 115074 800
rect 116122 0 116178 800
rect 117134 0 117190 800
rect 118238 0 118294 800
rect 119342 0 119398 800
rect 120446 0 120502 800
rect 121458 0 121514 800
rect 122562 0 122618 800
rect 123666 0 123722 800
rect 124770 0 124826 800
rect 125782 0 125838 800
rect 126886 0 126942 800
rect 127990 0 128046 800
rect 129094 0 129150 800
rect 130106 0 130162 800
rect 131210 0 131266 800
rect 132314 0 132370 800
rect 133418 0 133474 800
rect 134430 0 134486 800
rect 135534 0 135590 800
rect 136638 0 136694 800
rect 137742 0 137798 800
rect 138754 0 138810 800
rect 139858 0 139914 800
rect 140962 0 141018 800
rect 142066 0 142122 800
rect 143078 0 143134 800
rect 144182 0 144238 800
rect 145286 0 145342 800
rect 146390 0 146446 800
rect 147402 0 147458 800
rect 148506 0 148562 800
rect 149610 0 149666 800
rect 150714 0 150770 800
rect 151726 0 151782 800
rect 152830 0 152886 800
rect 153934 0 153990 800
rect 155038 0 155094 800
rect 156050 0 156106 800
rect 157154 0 157210 800
rect 158258 0 158314 800
rect 159362 0 159418 800
rect 160374 0 160430 800
rect 161478 0 161534 800
rect 162582 0 162638 800
rect 163686 0 163742 800
rect 164698 0 164754 800
rect 165802 0 165858 800
rect 166906 0 166962 800
rect 168010 0 168066 800
rect 169022 0 169078 800
rect 170126 0 170182 800
rect 171230 0 171286 800
rect 172334 0 172390 800
rect 173346 0 173402 800
rect 174450 0 174506 800
rect 175554 0 175610 800
rect 176658 0 176714 800
rect 177670 0 177726 800
rect 178774 0 178830 800
rect 179878 0 179934 800
rect 180982 0 181038 800
rect 181994 0 182050 800
rect 183098 0 183154 800
rect 184202 0 184258 800
rect 185306 0 185362 800
rect 186318 0 186374 800
rect 187422 0 187478 800
rect 188526 0 188582 800
rect 189630 0 189686 800
rect 190642 0 190698 800
rect 191746 0 191802 800
rect 192850 0 192906 800
rect 193954 0 194010 800
rect 194966 0 195022 800
rect 196070 0 196126 800
rect 197174 0 197230 800
rect 198278 0 198334 800
rect 199290 0 199346 800
rect 200394 0 200450 800
rect 201498 0 201554 800
rect 202602 0 202658 800
rect 203614 0 203670 800
rect 204718 0 204774 800
rect 205822 0 205878 800
rect 206926 0 206982 800
rect 207938 0 207994 800
rect 209042 0 209098 800
rect 210146 0 210202 800
rect 211250 0 211306 800
rect 212262 0 212318 800
rect 213366 0 213422 800
rect 214470 0 214526 800
rect 215574 0 215630 800
rect 216586 0 216642 800
rect 217690 0 217746 800
rect 218794 0 218850 800
rect 219898 0 219954 800
rect 220910 0 220966 800
rect 222014 0 222070 800
rect 223118 0 223174 800
rect 224222 0 224278 800
rect 225234 0 225290 800
rect 226338 0 226394 800
rect 227442 0 227498 800
rect 228546 0 228602 800
rect 229558 0 229614 800
rect 230662 0 230718 800
rect 231766 0 231822 800
rect 232870 0 232926 800
rect 233882 0 233938 800
rect 234986 0 235042 800
rect 236090 0 236146 800
rect 237194 0 237250 800
rect 238206 0 238262 800
rect 239310 0 239366 800
rect 240414 0 240470 800
rect 241518 0 241574 800
rect 242530 0 242586 800
rect 243634 0 243690 800
rect 244738 0 244794 800
rect 245842 0 245898 800
rect 246854 0 246910 800
rect 247958 0 248014 800
rect 249062 0 249118 800
rect 250166 0 250222 800
rect 251178 0 251234 800
rect 252282 0 252338 800
rect 253386 0 253442 800
rect 254490 0 254546 800
rect 255502 0 255558 800
rect 256606 0 256662 800
rect 257710 0 257766 800
rect 258814 0 258870 800
rect 259826 0 259882 800
rect 260930 0 260986 800
rect 262034 0 262090 800
rect 263138 0 263194 800
rect 264150 0 264206 800
rect 265254 0 265310 800
rect 266358 0 266414 800
rect 267462 0 267518 800
rect 268474 0 268530 800
rect 269578 0 269634 800
rect 270682 0 270738 800
rect 271786 0 271842 800
rect 272798 0 272854 800
rect 273902 0 273958 800
rect 275006 0 275062 800
rect 276110 0 276166 800
rect 277122 0 277178 800
rect 278226 0 278282 800
rect 279330 0 279386 800
<< obsm2 >>
rect 20 856 279384 299849
rect 20 2 422 856
rect 590 2 1434 856
rect 1602 2 2538 856
rect 2706 2 3642 856
rect 3810 2 4654 856
rect 4822 2 5758 856
rect 5926 2 6862 856
rect 7030 2 7966 856
rect 8134 2 8978 856
rect 9146 2 10082 856
rect 10250 2 11186 856
rect 11354 2 12290 856
rect 12458 2 13302 856
rect 13470 2 14406 856
rect 14574 2 15510 856
rect 15678 2 16614 856
rect 16782 2 17626 856
rect 17794 2 18730 856
rect 18898 2 19834 856
rect 20002 2 20938 856
rect 21106 2 21950 856
rect 22118 2 23054 856
rect 23222 2 24158 856
rect 24326 2 25262 856
rect 25430 2 26274 856
rect 26442 2 27378 856
rect 27546 2 28482 856
rect 28650 2 29586 856
rect 29754 2 30598 856
rect 30766 2 31702 856
rect 31870 2 32806 856
rect 32974 2 33910 856
rect 34078 2 34922 856
rect 35090 2 36026 856
rect 36194 2 37130 856
rect 37298 2 38234 856
rect 38402 2 39246 856
rect 39414 2 40350 856
rect 40518 2 41454 856
rect 41622 2 42558 856
rect 42726 2 43570 856
rect 43738 2 44674 856
rect 44842 2 45778 856
rect 45946 2 46882 856
rect 47050 2 47894 856
rect 48062 2 48998 856
rect 49166 2 50102 856
rect 50270 2 51206 856
rect 51374 2 52218 856
rect 52386 2 53322 856
rect 53490 2 54426 856
rect 54594 2 55530 856
rect 55698 2 56542 856
rect 56710 2 57646 856
rect 57814 2 58750 856
rect 58918 2 59854 856
rect 60022 2 60866 856
rect 61034 2 61970 856
rect 62138 2 63074 856
rect 63242 2 64178 856
rect 64346 2 65190 856
rect 65358 2 66294 856
rect 66462 2 67398 856
rect 67566 2 68502 856
rect 68670 2 69514 856
rect 69682 2 70618 856
rect 70786 2 71722 856
rect 71890 2 72826 856
rect 72994 2 73838 856
rect 74006 2 74942 856
rect 75110 2 76046 856
rect 76214 2 77150 856
rect 77318 2 78162 856
rect 78330 2 79266 856
rect 79434 2 80370 856
rect 80538 2 81474 856
rect 81642 2 82486 856
rect 82654 2 83590 856
rect 83758 2 84694 856
rect 84862 2 85798 856
rect 85966 2 86810 856
rect 86978 2 87914 856
rect 88082 2 89018 856
rect 89186 2 90122 856
rect 90290 2 91134 856
rect 91302 2 92238 856
rect 92406 2 93342 856
rect 93510 2 94446 856
rect 94614 2 95458 856
rect 95626 2 96562 856
rect 96730 2 97666 856
rect 97834 2 98770 856
rect 98938 2 99782 856
rect 99950 2 100886 856
rect 101054 2 101990 856
rect 102158 2 103094 856
rect 103262 2 104106 856
rect 104274 2 105210 856
rect 105378 2 106314 856
rect 106482 2 107418 856
rect 107586 2 108430 856
rect 108598 2 109534 856
rect 109702 2 110638 856
rect 110806 2 111742 856
rect 111910 2 112754 856
rect 112922 2 113858 856
rect 114026 2 114962 856
rect 115130 2 116066 856
rect 116234 2 117078 856
rect 117246 2 118182 856
rect 118350 2 119286 856
rect 119454 2 120390 856
rect 120558 2 121402 856
rect 121570 2 122506 856
rect 122674 2 123610 856
rect 123778 2 124714 856
rect 124882 2 125726 856
rect 125894 2 126830 856
rect 126998 2 127934 856
rect 128102 2 129038 856
rect 129206 2 130050 856
rect 130218 2 131154 856
rect 131322 2 132258 856
rect 132426 2 133362 856
rect 133530 2 134374 856
rect 134542 2 135478 856
rect 135646 2 136582 856
rect 136750 2 137686 856
rect 137854 2 138698 856
rect 138866 2 139802 856
rect 139970 2 140906 856
rect 141074 2 142010 856
rect 142178 2 143022 856
rect 143190 2 144126 856
rect 144294 2 145230 856
rect 145398 2 146334 856
rect 146502 2 147346 856
rect 147514 2 148450 856
rect 148618 2 149554 856
rect 149722 2 150658 856
rect 150826 2 151670 856
rect 151838 2 152774 856
rect 152942 2 153878 856
rect 154046 2 154982 856
rect 155150 2 155994 856
rect 156162 2 157098 856
rect 157266 2 158202 856
rect 158370 2 159306 856
rect 159474 2 160318 856
rect 160486 2 161422 856
rect 161590 2 162526 856
rect 162694 2 163630 856
rect 163798 2 164642 856
rect 164810 2 165746 856
rect 165914 2 166850 856
rect 167018 2 167954 856
rect 168122 2 168966 856
rect 169134 2 170070 856
rect 170238 2 171174 856
rect 171342 2 172278 856
rect 172446 2 173290 856
rect 173458 2 174394 856
rect 174562 2 175498 856
rect 175666 2 176602 856
rect 176770 2 177614 856
rect 177782 2 178718 856
rect 178886 2 179822 856
rect 179990 2 180926 856
rect 181094 2 181938 856
rect 182106 2 183042 856
rect 183210 2 184146 856
rect 184314 2 185250 856
rect 185418 2 186262 856
rect 186430 2 187366 856
rect 187534 2 188470 856
rect 188638 2 189574 856
rect 189742 2 190586 856
rect 190754 2 191690 856
rect 191858 2 192794 856
rect 192962 2 193898 856
rect 194066 2 194910 856
rect 195078 2 196014 856
rect 196182 2 197118 856
rect 197286 2 198222 856
rect 198390 2 199234 856
rect 199402 2 200338 856
rect 200506 2 201442 856
rect 201610 2 202546 856
rect 202714 2 203558 856
rect 203726 2 204662 856
rect 204830 2 205766 856
rect 205934 2 206870 856
rect 207038 2 207882 856
rect 208050 2 208986 856
rect 209154 2 210090 856
rect 210258 2 211194 856
rect 211362 2 212206 856
rect 212374 2 213310 856
rect 213478 2 214414 856
rect 214582 2 215518 856
rect 215686 2 216530 856
rect 216698 2 217634 856
rect 217802 2 218738 856
rect 218906 2 219842 856
rect 220010 2 220854 856
rect 221022 2 221958 856
rect 222126 2 223062 856
rect 223230 2 224166 856
rect 224334 2 225178 856
rect 225346 2 226282 856
rect 226450 2 227386 856
rect 227554 2 228490 856
rect 228658 2 229502 856
rect 229670 2 230606 856
rect 230774 2 231710 856
rect 231878 2 232814 856
rect 232982 2 233826 856
rect 233994 2 234930 856
rect 235098 2 236034 856
rect 236202 2 237138 856
rect 237306 2 238150 856
rect 238318 2 239254 856
rect 239422 2 240358 856
rect 240526 2 241462 856
rect 241630 2 242474 856
rect 242642 2 243578 856
rect 243746 2 244682 856
rect 244850 2 245786 856
rect 245954 2 246798 856
rect 246966 2 247902 856
rect 248070 2 249006 856
rect 249174 2 250110 856
rect 250278 2 251122 856
rect 251290 2 252226 856
rect 252394 2 253330 856
rect 253498 2 254434 856
rect 254602 2 255446 856
rect 255614 2 256550 856
rect 256718 2 257654 856
rect 257822 2 258758 856
rect 258926 2 259770 856
rect 259938 2 260874 856
rect 261042 2 261978 856
rect 262146 2 263082 856
rect 263250 2 264094 856
rect 264262 2 265198 856
rect 265366 2 266302 856
rect 266470 2 267406 856
rect 267574 2 268418 856
rect 268586 2 269522 856
rect 269690 2 270626 856
rect 270794 2 271730 856
rect 271898 2 272742 856
rect 272910 2 273846 856
rect 274014 2 274950 856
rect 275118 2 276054 856
rect 276222 2 277066 856
rect 277234 2 278170 856
rect 278338 2 279274 856
<< metal3 >>
rect 0 299752 800 299872
rect 0 299344 800 299464
rect 0 299072 800 299192
rect 0 298664 800 298784
rect 0 298256 800 298376
rect 0 297984 800 298104
rect 0 297576 800 297696
rect 0 297168 800 297288
rect 0 296896 800 297016
rect 0 296488 800 296608
rect 0 296216 800 296336
rect 0 295808 800 295928
rect 0 295400 800 295520
rect 0 295128 800 295248
rect 0 294720 800 294840
rect 0 294312 800 294432
rect 0 294040 800 294160
rect 0 293632 800 293752
rect 0 293360 800 293480
rect 0 292952 800 293072
rect 0 292544 800 292664
rect 0 292272 800 292392
rect 0 291864 800 291984
rect 0 291456 800 291576
rect 0 291184 800 291304
rect 0 290776 800 290896
rect 0 290504 800 290624
rect 0 290096 800 290216
rect 0 289688 800 289808
rect 0 289416 800 289536
rect 0 289008 800 289128
rect 0 288600 800 288720
rect 0 288328 800 288448
rect 0 287920 800 288040
rect 0 287648 800 287768
rect 0 287240 800 287360
rect 0 286832 800 286952
rect 0 286560 800 286680
rect 0 286152 800 286272
rect 0 285744 800 285864
rect 0 285472 800 285592
rect 0 285064 800 285184
rect 0 284792 800 284912
rect 0 284384 800 284504
rect 0 283976 800 284096
rect 0 283704 800 283824
rect 0 283296 800 283416
rect 0 282888 800 283008
rect 0 282616 800 282736
rect 0 282208 800 282328
rect 0 281936 800 282056
rect 0 281528 800 281648
rect 0 281120 800 281240
rect 0 280848 800 280968
rect 0 280440 800 280560
rect 0 280032 800 280152
rect 0 279760 800 279880
rect 0 279352 800 279472
rect 0 279080 800 279200
rect 0 278672 800 278792
rect 0 278264 800 278384
rect 0 277992 800 278112
rect 0 277584 800 277704
rect 0 277176 800 277296
rect 0 276904 800 277024
rect 0 276496 800 276616
rect 0 276224 800 276344
rect 0 275816 800 275936
rect 0 275408 800 275528
rect 0 275136 800 275256
rect 0 274728 800 274848
rect 0 274320 800 274440
rect 0 274048 800 274168
rect 0 273640 800 273760
rect 0 273368 800 273488
rect 0 272960 800 273080
rect 0 272552 800 272672
rect 0 272280 800 272400
rect 0 271872 800 271992
rect 0 271464 800 271584
rect 0 271192 800 271312
rect 0 270784 800 270904
rect 0 270512 800 270632
rect 0 270104 800 270224
rect 0 269696 800 269816
rect 0 269424 800 269544
rect 0 269016 800 269136
rect 0 268608 800 268728
rect 0 268336 800 268456
rect 0 267928 800 268048
rect 0 267656 800 267776
rect 0 267248 800 267368
rect 0 266840 800 266960
rect 0 266568 800 266688
rect 0 266160 800 266280
rect 0 265752 800 265872
rect 0 265480 800 265600
rect 0 265072 800 265192
rect 0 264800 800 264920
rect 0 264392 800 264512
rect 0 263984 800 264104
rect 0 263712 800 263832
rect 0 263304 800 263424
rect 0 262896 800 263016
rect 0 262624 800 262744
rect 0 262216 800 262336
rect 0 261808 800 261928
rect 0 261536 800 261656
rect 0 261128 800 261248
rect 0 260856 800 260976
rect 0 260448 800 260568
rect 0 260040 800 260160
rect 0 259768 800 259888
rect 0 259360 800 259480
rect 0 258952 800 259072
rect 0 258680 800 258800
rect 0 258272 800 258392
rect 0 258000 800 258120
rect 0 257592 800 257712
rect 0 257184 800 257304
rect 0 256912 800 257032
rect 0 256504 800 256624
rect 0 256096 800 256216
rect 0 255824 800 255944
rect 0 255416 800 255536
rect 0 255144 800 255264
rect 0 254736 800 254856
rect 0 254328 800 254448
rect 0 254056 800 254176
rect 0 253648 800 253768
rect 0 253240 800 253360
rect 0 252968 800 253088
rect 0 252560 800 252680
rect 0 252288 800 252408
rect 0 251880 800 252000
rect 0 251472 800 251592
rect 0 251200 800 251320
rect 0 250792 800 250912
rect 0 250384 800 250504
rect 0 250112 800 250232
rect 0 249704 800 249824
rect 0 249432 800 249552
rect 0 249024 800 249144
rect 0 248616 800 248736
rect 0 248344 800 248464
rect 0 247936 800 248056
rect 0 247528 800 247648
rect 0 247256 800 247376
rect 0 246848 800 246968
rect 0 246576 800 246696
rect 0 246168 800 246288
rect 0 245760 800 245880
rect 0 245488 800 245608
rect 0 245080 800 245200
rect 0 244672 800 244792
rect 0 244400 800 244520
rect 0 243992 800 244112
rect 0 243720 800 243840
rect 0 243312 800 243432
rect 0 242904 800 243024
rect 0 242632 800 242752
rect 0 242224 800 242344
rect 0 241816 800 241936
rect 0 241544 800 241664
rect 0 241136 800 241256
rect 0 240864 800 240984
rect 0 240456 800 240576
rect 0 240048 800 240168
rect 0 239776 800 239896
rect 0 239368 800 239488
rect 0 238960 800 239080
rect 0 238688 800 238808
rect 0 238280 800 238400
rect 0 238008 800 238128
rect 0 237600 800 237720
rect 0 237192 800 237312
rect 0 236920 800 237040
rect 0 236512 800 236632
rect 0 236104 800 236224
rect 0 235832 800 235952
rect 0 235424 800 235544
rect 0 235152 800 235272
rect 0 234744 800 234864
rect 0 234336 800 234456
rect 0 234064 800 234184
rect 0 233656 800 233776
rect 0 233248 800 233368
rect 0 232976 800 233096
rect 0 232568 800 232688
rect 0 232296 800 232416
rect 0 231888 800 232008
rect 0 231480 800 231600
rect 0 231208 800 231328
rect 0 230800 800 230920
rect 0 230392 800 230512
rect 0 230120 800 230240
rect 0 229712 800 229832
rect 0 229440 800 229560
rect 0 229032 800 229152
rect 0 228624 800 228744
rect 0 228352 800 228472
rect 0 227944 800 228064
rect 0 227536 800 227656
rect 0 227264 800 227384
rect 0 226856 800 226976
rect 0 226584 800 226704
rect 0 226176 800 226296
rect 0 225768 800 225888
rect 0 225496 800 225616
rect 0 225088 800 225208
rect 0 224680 800 224800
rect 0 224408 800 224528
rect 0 224000 800 224120
rect 0 223592 800 223712
rect 0 223320 800 223440
rect 0 222912 800 223032
rect 0 222640 800 222760
rect 0 222232 800 222352
rect 0 221824 800 221944
rect 0 221552 800 221672
rect 0 221144 800 221264
rect 0 220736 800 220856
rect 0 220464 800 220584
rect 0 220056 800 220176
rect 0 219784 800 219904
rect 0 219376 800 219496
rect 0 218968 800 219088
rect 0 218696 800 218816
rect 0 218288 800 218408
rect 0 217880 800 218000
rect 0 217608 800 217728
rect 0 217200 800 217320
rect 0 216928 800 217048
rect 0 216520 800 216640
rect 0 216112 800 216232
rect 0 215840 800 215960
rect 0 215432 800 215552
rect 0 215024 800 215144
rect 0 214752 800 214872
rect 0 214344 800 214464
rect 0 214072 800 214192
rect 0 213664 800 213784
rect 0 213256 800 213376
rect 0 212984 800 213104
rect 0 212576 800 212696
rect 0 212168 800 212288
rect 0 211896 800 212016
rect 0 211488 800 211608
rect 0 211216 800 211336
rect 0 210808 800 210928
rect 0 210400 800 210520
rect 0 210128 800 210248
rect 0 209720 800 209840
rect 0 209312 800 209432
rect 0 209040 800 209160
rect 0 208632 800 208752
rect 0 208360 800 208480
rect 0 207952 800 208072
rect 0 207544 800 207664
rect 0 207272 800 207392
rect 0 206864 800 206984
rect 0 206456 800 206576
rect 0 206184 800 206304
rect 0 205776 800 205896
rect 0 205504 800 205624
rect 0 205096 800 205216
rect 0 204688 800 204808
rect 0 204416 800 204536
rect 0 204008 800 204128
rect 0 203600 800 203720
rect 0 203328 800 203448
rect 0 202920 800 203040
rect 0 202648 800 202768
rect 0 202240 800 202360
rect 0 201832 800 201952
rect 0 201560 800 201680
rect 0 201152 800 201272
rect 0 200744 800 200864
rect 0 200472 800 200592
rect 0 200064 800 200184
rect 0 199792 800 199912
rect 0 199384 800 199504
rect 0 198976 800 199096
rect 0 198704 800 198824
rect 0 198296 800 198416
rect 0 197888 800 198008
rect 0 197616 800 197736
rect 0 197208 800 197328
rect 0 196936 800 197056
rect 0 196528 800 196648
rect 0 196120 800 196240
rect 0 195848 800 195968
rect 0 195440 800 195560
rect 0 195032 800 195152
rect 0 194760 800 194880
rect 0 194352 800 194472
rect 0 194080 800 194200
rect 0 193672 800 193792
rect 0 193264 800 193384
rect 0 192992 800 193112
rect 0 192584 800 192704
rect 0 192176 800 192296
rect 0 191904 800 192024
rect 0 191496 800 191616
rect 0 191224 800 191344
rect 0 190816 800 190936
rect 0 190408 800 190528
rect 0 190136 800 190256
rect 0 189728 800 189848
rect 0 189320 800 189440
rect 0 189048 800 189168
rect 0 188640 800 188760
rect 0 188368 800 188488
rect 0 187960 800 188080
rect 0 187552 800 187672
rect 0 187280 800 187400
rect 0 186872 800 186992
rect 0 186464 800 186584
rect 0 186192 800 186312
rect 0 185784 800 185904
rect 0 185376 800 185496
rect 0 185104 800 185224
rect 0 184696 800 184816
rect 0 184424 800 184544
rect 0 184016 800 184136
rect 0 183608 800 183728
rect 0 183336 800 183456
rect 0 182928 800 183048
rect 0 182520 800 182640
rect 0 182248 800 182368
rect 0 181840 800 181960
rect 0 181568 800 181688
rect 0 181160 800 181280
rect 0 180752 800 180872
rect 0 180480 800 180600
rect 0 180072 800 180192
rect 0 179664 800 179784
rect 0 179392 800 179512
rect 0 178984 800 179104
rect 0 178712 800 178832
rect 0 178304 800 178424
rect 0 177896 800 178016
rect 0 177624 800 177744
rect 0 177216 800 177336
rect 0 176808 800 176928
rect 0 176536 800 176656
rect 0 176128 800 176248
rect 0 175856 800 175976
rect 0 175448 800 175568
rect 0 175040 800 175160
rect 0 174768 800 174888
rect 0 174360 800 174480
rect 0 173952 800 174072
rect 0 173680 800 173800
rect 0 173272 800 173392
rect 0 173000 800 173120
rect 0 172592 800 172712
rect 0 172184 800 172304
rect 0 171912 800 172032
rect 0 171504 800 171624
rect 0 171096 800 171216
rect 0 170824 800 170944
rect 0 170416 800 170536
rect 0 170144 800 170264
rect 0 169736 800 169856
rect 0 169328 800 169448
rect 0 169056 800 169176
rect 0 168648 800 168768
rect 0 168240 800 168360
rect 0 167968 800 168088
rect 0 167560 800 167680
rect 0 167288 800 167408
rect 0 166880 800 167000
rect 0 166472 800 166592
rect 0 166200 800 166320
rect 0 165792 800 165912
rect 0 165384 800 165504
rect 0 165112 800 165232
rect 0 164704 800 164824
rect 0 164432 800 164552
rect 0 164024 800 164144
rect 0 163616 800 163736
rect 0 163344 800 163464
rect 0 162936 800 163056
rect 0 162528 800 162648
rect 0 162256 800 162376
rect 0 161848 800 161968
rect 0 161576 800 161696
rect 0 161168 800 161288
rect 0 160760 800 160880
rect 0 160488 800 160608
rect 0 160080 800 160200
rect 0 159672 800 159792
rect 0 159400 800 159520
rect 0 158992 800 159112
rect 0 158720 800 158840
rect 0 158312 800 158432
rect 0 157904 800 158024
rect 0 157632 800 157752
rect 0 157224 800 157344
rect 0 156816 800 156936
rect 0 156544 800 156664
rect 0 156136 800 156256
rect 0 155864 800 155984
rect 0 155456 800 155576
rect 0 155048 800 155168
rect 0 154776 800 154896
rect 0 154368 800 154488
rect 0 153960 800 154080
rect 0 153688 800 153808
rect 0 153280 800 153400
rect 0 153008 800 153128
rect 0 152600 800 152720
rect 0 152192 800 152312
rect 0 151920 800 152040
rect 0 151512 800 151632
rect 0 151104 800 151224
rect 0 150832 800 150952
rect 0 150424 800 150544
rect 0 150152 800 150272
rect 0 149744 800 149864
rect 0 149336 800 149456
rect 0 149064 800 149184
rect 0 148656 800 148776
rect 0 148248 800 148368
rect 0 147976 800 148096
rect 0 147568 800 147688
rect 0 147160 800 147280
rect 0 146888 800 147008
rect 0 146480 800 146600
rect 0 146208 800 146328
rect 0 145800 800 145920
rect 0 145392 800 145512
rect 0 145120 800 145240
rect 0 144712 800 144832
rect 0 144304 800 144424
rect 0 144032 800 144152
rect 0 143624 800 143744
rect 0 143352 800 143472
rect 0 142944 800 143064
rect 0 142536 800 142656
rect 0 142264 800 142384
rect 0 141856 800 141976
rect 0 141448 800 141568
rect 0 141176 800 141296
rect 0 140768 800 140888
rect 0 140496 800 140616
rect 0 140088 800 140208
rect 0 139680 800 139800
rect 0 139408 800 139528
rect 0 139000 800 139120
rect 0 138592 800 138712
rect 0 138320 800 138440
rect 0 137912 800 138032
rect 0 137640 800 137760
rect 0 137232 800 137352
rect 0 136824 800 136944
rect 0 136552 800 136672
rect 0 136144 800 136264
rect 0 135736 800 135856
rect 0 135464 800 135584
rect 0 135056 800 135176
rect 0 134784 800 134904
rect 0 134376 800 134496
rect 0 133968 800 134088
rect 0 133696 800 133816
rect 0 133288 800 133408
rect 0 132880 800 133000
rect 0 132608 800 132728
rect 0 132200 800 132320
rect 0 131928 800 132048
rect 0 131520 800 131640
rect 0 131112 800 131232
rect 0 130840 800 130960
rect 0 130432 800 130552
rect 0 130024 800 130144
rect 0 129752 800 129872
rect 0 129344 800 129464
rect 0 129072 800 129192
rect 0 128664 800 128784
rect 0 128256 800 128376
rect 0 127984 800 128104
rect 0 127576 800 127696
rect 0 127168 800 127288
rect 0 126896 800 127016
rect 0 126488 800 126608
rect 0 126216 800 126336
rect 0 125808 800 125928
rect 0 125400 800 125520
rect 0 125128 800 125248
rect 0 124720 800 124840
rect 0 124312 800 124432
rect 0 124040 800 124160
rect 0 123632 800 123752
rect 0 123360 800 123480
rect 0 122952 800 123072
rect 0 122544 800 122664
rect 0 122272 800 122392
rect 0 121864 800 121984
rect 0 121456 800 121576
rect 0 121184 800 121304
rect 0 120776 800 120896
rect 0 120504 800 120624
rect 0 120096 800 120216
rect 0 119688 800 119808
rect 0 119416 800 119536
rect 0 119008 800 119128
rect 0 118600 800 118720
rect 0 118328 800 118448
rect 0 117920 800 118040
rect 0 117648 800 117768
rect 0 117240 800 117360
rect 0 116832 800 116952
rect 0 116560 800 116680
rect 0 116152 800 116272
rect 0 115744 800 115864
rect 0 115472 800 115592
rect 0 115064 800 115184
rect 0 114792 800 114912
rect 0 114384 800 114504
rect 0 113976 800 114096
rect 0 113704 800 113824
rect 0 113296 800 113416
rect 0 112888 800 113008
rect 0 112616 800 112736
rect 0 112208 800 112328
rect 0 111800 800 111920
rect 0 111528 800 111648
rect 0 111120 800 111240
rect 0 110848 800 110968
rect 0 110440 800 110560
rect 0 110032 800 110152
rect 0 109760 800 109880
rect 0 109352 800 109472
rect 0 108944 800 109064
rect 0 108672 800 108792
rect 0 108264 800 108384
rect 0 107992 800 108112
rect 0 107584 800 107704
rect 0 107176 800 107296
rect 0 106904 800 107024
rect 0 106496 800 106616
rect 0 106088 800 106208
rect 0 105816 800 105936
rect 0 105408 800 105528
rect 0 105136 800 105256
rect 0 104728 800 104848
rect 0 104320 800 104440
rect 0 104048 800 104168
rect 0 103640 800 103760
rect 0 103232 800 103352
rect 0 102960 800 103080
rect 0 102552 800 102672
rect 0 102280 800 102400
rect 0 101872 800 101992
rect 0 101464 800 101584
rect 0 101192 800 101312
rect 0 100784 800 100904
rect 0 100376 800 100496
rect 0 100104 800 100224
rect 0 99696 800 99816
rect 0 99424 800 99544
rect 0 99016 800 99136
rect 0 98608 800 98728
rect 0 98336 800 98456
rect 0 97928 800 98048
rect 0 97520 800 97640
rect 0 97248 800 97368
rect 0 96840 800 96960
rect 0 96568 800 96688
rect 0 96160 800 96280
rect 0 95752 800 95872
rect 0 95480 800 95600
rect 0 95072 800 95192
rect 0 94664 800 94784
rect 0 94392 800 94512
rect 0 93984 800 94104
rect 0 93712 800 93832
rect 0 93304 800 93424
rect 0 92896 800 93016
rect 0 92624 800 92744
rect 0 92216 800 92336
rect 0 91808 800 91928
rect 0 91536 800 91656
rect 0 91128 800 91248
rect 0 90856 800 90976
rect 0 90448 800 90568
rect 0 90040 800 90160
rect 0 89768 800 89888
rect 0 89360 800 89480
rect 0 88952 800 89072
rect 0 88680 800 88800
rect 0 88272 800 88392
rect 0 88000 800 88120
rect 0 87592 800 87712
rect 0 87184 800 87304
rect 0 86912 800 87032
rect 0 86504 800 86624
rect 0 86096 800 86216
rect 0 85824 800 85944
rect 0 85416 800 85536
rect 0 85144 800 85264
rect 0 84736 800 84856
rect 0 84328 800 84448
rect 0 84056 800 84176
rect 0 83648 800 83768
rect 0 83240 800 83360
rect 0 82968 800 83088
rect 0 82560 800 82680
rect 0 82288 800 82408
rect 0 81880 800 82000
rect 0 81472 800 81592
rect 0 81200 800 81320
rect 0 80792 800 80912
rect 0 80384 800 80504
rect 0 80112 800 80232
rect 0 79704 800 79824
rect 0 79432 800 79552
rect 0 79024 800 79144
rect 0 78616 800 78736
rect 0 78344 800 78464
rect 0 77936 800 78056
rect 0 77528 800 77648
rect 0 77256 800 77376
rect 0 76848 800 76968
rect 0 76576 800 76696
rect 0 76168 800 76288
rect 0 75760 800 75880
rect 0 75488 800 75608
rect 0 75080 800 75200
rect 0 74672 800 74792
rect 0 74400 800 74520
rect 0 73992 800 74112
rect 0 73584 800 73704
rect 0 73312 800 73432
rect 0 72904 800 73024
rect 0 72632 800 72752
rect 0 72224 800 72344
rect 0 71816 800 71936
rect 0 71544 800 71664
rect 0 71136 800 71256
rect 0 70728 800 70848
rect 0 70456 800 70576
rect 0 70048 800 70168
rect 0 69776 800 69896
rect 0 69368 800 69488
rect 0 68960 800 69080
rect 0 68688 800 68808
rect 0 68280 800 68400
rect 0 67872 800 67992
rect 0 67600 800 67720
rect 0 67192 800 67312
rect 0 66920 800 67040
rect 0 66512 800 66632
rect 0 66104 800 66224
rect 0 65832 800 65952
rect 0 65424 800 65544
rect 0 65016 800 65136
rect 0 64744 800 64864
rect 0 64336 800 64456
rect 0 64064 800 64184
rect 0 63656 800 63776
rect 0 63248 800 63368
rect 0 62976 800 63096
rect 0 62568 800 62688
rect 0 62160 800 62280
rect 0 61888 800 62008
rect 0 61480 800 61600
rect 0 61208 800 61328
rect 0 60800 800 60920
rect 0 60392 800 60512
rect 0 60120 800 60240
rect 0 59712 800 59832
rect 0 59304 800 59424
rect 0 59032 800 59152
rect 0 58624 800 58744
rect 0 58352 800 58472
rect 0 57944 800 58064
rect 0 57536 800 57656
rect 0 57264 800 57384
rect 0 56856 800 56976
rect 0 56448 800 56568
rect 0 56176 800 56296
rect 0 55768 800 55888
rect 0 55496 800 55616
rect 0 55088 800 55208
rect 0 54680 800 54800
rect 0 54408 800 54528
rect 0 54000 800 54120
rect 0 53592 800 53712
rect 0 53320 800 53440
rect 0 52912 800 53032
rect 0 52640 800 52760
rect 0 52232 800 52352
rect 0 51824 800 51944
rect 0 51552 800 51672
rect 0 51144 800 51264
rect 0 50736 800 50856
rect 0 50464 800 50584
rect 0 50056 800 50176
rect 0 49784 800 49904
rect 0 49376 800 49496
rect 0 48968 800 49088
rect 0 48696 800 48816
rect 0 48288 800 48408
rect 0 47880 800 48000
rect 0 47608 800 47728
rect 0 47200 800 47320
rect 0 46928 800 47048
rect 0 46520 800 46640
rect 0 46112 800 46232
rect 0 45840 800 45960
rect 0 45432 800 45552
rect 0 45024 800 45144
rect 0 44752 800 44872
rect 0 44344 800 44464
rect 0 44072 800 44192
rect 0 43664 800 43784
rect 0 43256 800 43376
rect 0 42984 800 43104
rect 0 42576 800 42696
rect 0 42168 800 42288
rect 0 41896 800 42016
rect 0 41488 800 41608
rect 0 41216 800 41336
rect 0 40808 800 40928
rect 0 40400 800 40520
rect 0 40128 800 40248
rect 0 39720 800 39840
rect 0 39312 800 39432
rect 0 39040 800 39160
rect 0 38632 800 38752
rect 0 38360 800 38480
rect 0 37952 800 38072
rect 0 37544 800 37664
rect 0 37272 800 37392
rect 0 36864 800 36984
rect 0 36456 800 36576
rect 0 36184 800 36304
rect 0 35776 800 35896
rect 0 35368 800 35488
rect 0 35096 800 35216
rect 0 34688 800 34808
rect 0 34416 800 34536
rect 0 34008 800 34128
rect 0 33600 800 33720
rect 0 33328 800 33448
rect 0 32920 800 33040
rect 0 32512 800 32632
rect 0 32240 800 32360
rect 0 31832 800 31952
rect 0 31560 800 31680
rect 0 31152 800 31272
rect 0 30744 800 30864
rect 0 30472 800 30592
rect 0 30064 800 30184
rect 0 29656 800 29776
rect 0 29384 800 29504
rect 0 28976 800 29096
rect 0 28704 800 28824
rect 0 28296 800 28416
rect 0 27888 800 28008
rect 0 27616 800 27736
rect 0 27208 800 27328
rect 0 26800 800 26920
rect 0 26528 800 26648
rect 0 26120 800 26240
rect 0 25848 800 25968
rect 0 25440 800 25560
rect 0 25032 800 25152
rect 0 24760 800 24880
rect 0 24352 800 24472
rect 0 23944 800 24064
rect 0 23672 800 23792
rect 0 23264 800 23384
rect 0 22992 800 23112
rect 0 22584 800 22704
rect 0 22176 800 22296
rect 0 21904 800 22024
rect 0 21496 800 21616
rect 0 21088 800 21208
rect 0 20816 800 20936
rect 0 20408 800 20528
rect 0 20136 800 20256
rect 0 19728 800 19848
rect 0 19320 800 19440
rect 0 19048 800 19168
rect 0 18640 800 18760
rect 0 18232 800 18352
rect 0 17960 800 18080
rect 0 17552 800 17672
rect 0 17280 800 17400
rect 0 16872 800 16992
rect 0 16464 800 16584
rect 0 16192 800 16312
rect 0 15784 800 15904
rect 0 15376 800 15496
rect 0 15104 800 15224
rect 0 14696 800 14816
rect 0 14424 800 14544
rect 0 14016 800 14136
rect 0 13608 800 13728
rect 0 13336 800 13456
rect 0 12928 800 13048
rect 0 12520 800 12640
rect 0 12248 800 12368
rect 0 11840 800 11960
rect 0 11568 800 11688
rect 0 11160 800 11280
rect 0 10752 800 10872
rect 0 10480 800 10600
rect 0 10072 800 10192
rect 0 9664 800 9784
rect 0 9392 800 9512
rect 0 8984 800 9104
rect 0 8712 800 8832
rect 0 8304 800 8424
rect 0 7896 800 8016
rect 0 7624 800 7744
rect 0 7216 800 7336
rect 0 6808 800 6928
rect 0 6536 800 6656
rect 0 6128 800 6248
rect 0 5856 800 5976
rect 0 5448 800 5568
rect 0 5040 800 5160
rect 0 4768 800 4888
rect 0 4360 800 4480
rect 0 3952 800 4072
rect 0 3680 800 3800
rect 0 3272 800 3392
rect 0 3000 800 3120
rect 0 2592 800 2712
rect 0 2184 800 2304
rect 0 1912 800 2032
rect 0 1504 800 1624
rect 0 1096 800 1216
rect 0 824 800 944
rect 0 416 800 536
rect 0 144 800 264
<< obsm3 >>
rect 880 299672 275435 299845
rect 54 299544 275435 299672
rect 880 298992 275435 299544
rect 54 298864 275435 298992
rect 880 298584 275435 298864
rect 54 298456 275435 298584
rect 880 297904 275435 298456
rect 54 297776 275435 297904
rect 880 297496 275435 297776
rect 54 297368 275435 297496
rect 880 296816 275435 297368
rect 54 296688 275435 296816
rect 880 296136 275435 296688
rect 54 296008 275435 296136
rect 880 295728 275435 296008
rect 54 295600 275435 295728
rect 880 295048 275435 295600
rect 54 294920 275435 295048
rect 880 294640 275435 294920
rect 54 294512 275435 294640
rect 880 293960 275435 294512
rect 54 293832 275435 293960
rect 880 293280 275435 293832
rect 54 293152 275435 293280
rect 880 292872 275435 293152
rect 54 292744 275435 292872
rect 880 292192 275435 292744
rect 54 292064 275435 292192
rect 880 291784 275435 292064
rect 54 291656 275435 291784
rect 880 291104 275435 291656
rect 54 290976 275435 291104
rect 880 290424 275435 290976
rect 54 290296 275435 290424
rect 880 290016 275435 290296
rect 54 289888 275435 290016
rect 880 289336 275435 289888
rect 54 289208 275435 289336
rect 880 288928 275435 289208
rect 54 288800 275435 288928
rect 880 288248 275435 288800
rect 54 288120 275435 288248
rect 880 287568 275435 288120
rect 54 287440 275435 287568
rect 880 287160 275435 287440
rect 54 287032 275435 287160
rect 880 286480 275435 287032
rect 54 286352 275435 286480
rect 880 286072 275435 286352
rect 54 285944 275435 286072
rect 880 285392 275435 285944
rect 54 285264 275435 285392
rect 880 284712 275435 285264
rect 54 284584 275435 284712
rect 880 284304 275435 284584
rect 54 284176 275435 284304
rect 880 283624 275435 284176
rect 54 283496 275435 283624
rect 880 283216 275435 283496
rect 54 283088 275435 283216
rect 880 282536 275435 283088
rect 54 282408 275435 282536
rect 880 281856 275435 282408
rect 54 281728 275435 281856
rect 880 281448 275435 281728
rect 54 281320 275435 281448
rect 880 280768 275435 281320
rect 54 280640 275435 280768
rect 880 280360 275435 280640
rect 54 280232 275435 280360
rect 880 279680 275435 280232
rect 54 279552 275435 279680
rect 880 279000 275435 279552
rect 54 278872 275435 279000
rect 880 278592 275435 278872
rect 54 278464 275435 278592
rect 880 277912 275435 278464
rect 54 277784 275435 277912
rect 880 277504 275435 277784
rect 54 277376 275435 277504
rect 880 276824 275435 277376
rect 54 276696 275435 276824
rect 880 276144 275435 276696
rect 54 276016 275435 276144
rect 880 275736 275435 276016
rect 54 275608 275435 275736
rect 880 275056 275435 275608
rect 54 274928 275435 275056
rect 880 274648 275435 274928
rect 54 274520 275435 274648
rect 880 273968 275435 274520
rect 54 273840 275435 273968
rect 880 273288 275435 273840
rect 54 273160 275435 273288
rect 880 272880 275435 273160
rect 54 272752 275435 272880
rect 880 272200 275435 272752
rect 54 272072 275435 272200
rect 880 271792 275435 272072
rect 54 271664 275435 271792
rect 880 271112 275435 271664
rect 54 270984 275435 271112
rect 880 270432 275435 270984
rect 54 270304 275435 270432
rect 880 270024 275435 270304
rect 54 269896 275435 270024
rect 880 269344 275435 269896
rect 54 269216 275435 269344
rect 880 268936 275435 269216
rect 54 268808 275435 268936
rect 880 268256 275435 268808
rect 54 268128 275435 268256
rect 880 267576 275435 268128
rect 54 267448 275435 267576
rect 880 267168 275435 267448
rect 54 267040 275435 267168
rect 880 266488 275435 267040
rect 54 266360 275435 266488
rect 880 266080 275435 266360
rect 54 265952 275435 266080
rect 880 265400 275435 265952
rect 54 265272 275435 265400
rect 880 264720 275435 265272
rect 54 264592 275435 264720
rect 880 264312 275435 264592
rect 54 264184 275435 264312
rect 880 263632 275435 264184
rect 54 263504 275435 263632
rect 880 263224 275435 263504
rect 54 263096 275435 263224
rect 880 262544 275435 263096
rect 54 262416 275435 262544
rect 880 262136 275435 262416
rect 54 262008 275435 262136
rect 880 261456 275435 262008
rect 54 261328 275435 261456
rect 880 260776 275435 261328
rect 54 260648 275435 260776
rect 880 260368 275435 260648
rect 54 260240 275435 260368
rect 880 259688 275435 260240
rect 54 259560 275435 259688
rect 880 259280 275435 259560
rect 54 259152 275435 259280
rect 880 258600 275435 259152
rect 54 258472 275435 258600
rect 880 257920 275435 258472
rect 54 257792 275435 257920
rect 880 257512 275435 257792
rect 54 257384 275435 257512
rect 880 256832 275435 257384
rect 54 256704 275435 256832
rect 880 256424 275435 256704
rect 54 256296 275435 256424
rect 880 255744 275435 256296
rect 54 255616 275435 255744
rect 880 255064 275435 255616
rect 54 254936 275435 255064
rect 880 254656 275435 254936
rect 54 254528 275435 254656
rect 880 253976 275435 254528
rect 54 253848 275435 253976
rect 880 253568 275435 253848
rect 54 253440 275435 253568
rect 880 252888 275435 253440
rect 54 252760 275435 252888
rect 880 252208 275435 252760
rect 54 252080 275435 252208
rect 880 251800 275435 252080
rect 54 251672 275435 251800
rect 880 251120 275435 251672
rect 54 250992 275435 251120
rect 880 250712 275435 250992
rect 54 250584 275435 250712
rect 880 250032 275435 250584
rect 54 249904 275435 250032
rect 880 249352 275435 249904
rect 54 249224 275435 249352
rect 880 248944 275435 249224
rect 54 248816 275435 248944
rect 880 248264 275435 248816
rect 54 248136 275435 248264
rect 880 247856 275435 248136
rect 54 247728 275435 247856
rect 880 247176 275435 247728
rect 54 247048 275435 247176
rect 880 246496 275435 247048
rect 54 246368 275435 246496
rect 880 246088 275435 246368
rect 54 245960 275435 246088
rect 880 245408 275435 245960
rect 54 245280 275435 245408
rect 880 245000 275435 245280
rect 54 244872 275435 245000
rect 880 244320 275435 244872
rect 54 244192 275435 244320
rect 880 243640 275435 244192
rect 54 243512 275435 243640
rect 880 243232 275435 243512
rect 54 243104 275435 243232
rect 880 242552 275435 243104
rect 54 242424 275435 242552
rect 880 242144 275435 242424
rect 54 242016 275435 242144
rect 880 241464 275435 242016
rect 54 241336 275435 241464
rect 880 240784 275435 241336
rect 54 240656 275435 240784
rect 880 240376 275435 240656
rect 54 240248 275435 240376
rect 880 239696 275435 240248
rect 54 239568 275435 239696
rect 880 239288 275435 239568
rect 54 239160 275435 239288
rect 880 238608 275435 239160
rect 54 238480 275435 238608
rect 880 237928 275435 238480
rect 54 237800 275435 237928
rect 880 237520 275435 237800
rect 54 237392 275435 237520
rect 880 236840 275435 237392
rect 54 236712 275435 236840
rect 880 236432 275435 236712
rect 54 236304 275435 236432
rect 880 235752 275435 236304
rect 54 235624 275435 235752
rect 880 235072 275435 235624
rect 54 234944 275435 235072
rect 880 234664 275435 234944
rect 54 234536 275435 234664
rect 880 233984 275435 234536
rect 54 233856 275435 233984
rect 880 233576 275435 233856
rect 54 233448 275435 233576
rect 880 232896 275435 233448
rect 54 232768 275435 232896
rect 880 232216 275435 232768
rect 54 232088 275435 232216
rect 880 231808 275435 232088
rect 54 231680 275435 231808
rect 880 231128 275435 231680
rect 54 231000 275435 231128
rect 880 230720 275435 231000
rect 54 230592 275435 230720
rect 880 230040 275435 230592
rect 54 229912 275435 230040
rect 880 229360 275435 229912
rect 54 229232 275435 229360
rect 880 228952 275435 229232
rect 54 228824 275435 228952
rect 880 228272 275435 228824
rect 54 228144 275435 228272
rect 880 227864 275435 228144
rect 54 227736 275435 227864
rect 880 227184 275435 227736
rect 54 227056 275435 227184
rect 880 226504 275435 227056
rect 54 226376 275435 226504
rect 880 226096 275435 226376
rect 54 225968 275435 226096
rect 880 225416 275435 225968
rect 54 225288 275435 225416
rect 880 225008 275435 225288
rect 54 224880 275435 225008
rect 880 224328 275435 224880
rect 54 224200 275435 224328
rect 880 223920 275435 224200
rect 54 223792 275435 223920
rect 880 223240 275435 223792
rect 54 223112 275435 223240
rect 880 222560 275435 223112
rect 54 222432 275435 222560
rect 880 222152 275435 222432
rect 54 222024 275435 222152
rect 880 221472 275435 222024
rect 54 221344 275435 221472
rect 880 221064 275435 221344
rect 54 220936 275435 221064
rect 880 220384 275435 220936
rect 54 220256 275435 220384
rect 880 219704 275435 220256
rect 54 219576 275435 219704
rect 880 219296 275435 219576
rect 54 219168 275435 219296
rect 880 218616 275435 219168
rect 54 218488 275435 218616
rect 880 218208 275435 218488
rect 54 218080 275435 218208
rect 880 217528 275435 218080
rect 54 217400 275435 217528
rect 880 216848 275435 217400
rect 54 216720 275435 216848
rect 880 216440 275435 216720
rect 54 216312 275435 216440
rect 880 215760 275435 216312
rect 54 215632 275435 215760
rect 880 215352 275435 215632
rect 54 215224 275435 215352
rect 880 214672 275435 215224
rect 54 214544 275435 214672
rect 880 213992 275435 214544
rect 54 213864 275435 213992
rect 880 213584 275435 213864
rect 54 213456 275435 213584
rect 880 212904 275435 213456
rect 54 212776 275435 212904
rect 880 212496 275435 212776
rect 54 212368 275435 212496
rect 880 211816 275435 212368
rect 54 211688 275435 211816
rect 880 211136 275435 211688
rect 54 211008 275435 211136
rect 880 210728 275435 211008
rect 54 210600 275435 210728
rect 880 210048 275435 210600
rect 54 209920 275435 210048
rect 880 209640 275435 209920
rect 54 209512 275435 209640
rect 880 208960 275435 209512
rect 54 208832 275435 208960
rect 880 208280 275435 208832
rect 54 208152 275435 208280
rect 880 207872 275435 208152
rect 54 207744 275435 207872
rect 880 207192 275435 207744
rect 54 207064 275435 207192
rect 880 206784 275435 207064
rect 54 206656 275435 206784
rect 880 206104 275435 206656
rect 54 205976 275435 206104
rect 880 205424 275435 205976
rect 54 205296 275435 205424
rect 880 205016 275435 205296
rect 54 204888 275435 205016
rect 880 204336 275435 204888
rect 54 204208 275435 204336
rect 880 203928 275435 204208
rect 54 203800 275435 203928
rect 880 203248 275435 203800
rect 54 203120 275435 203248
rect 880 202568 275435 203120
rect 54 202440 275435 202568
rect 880 202160 275435 202440
rect 54 202032 275435 202160
rect 880 201480 275435 202032
rect 54 201352 275435 201480
rect 880 201072 275435 201352
rect 54 200944 275435 201072
rect 880 200392 275435 200944
rect 54 200264 275435 200392
rect 880 199712 275435 200264
rect 54 199584 275435 199712
rect 880 199304 275435 199584
rect 54 199176 275435 199304
rect 880 198624 275435 199176
rect 54 198496 275435 198624
rect 880 198216 275435 198496
rect 54 198088 275435 198216
rect 880 197536 275435 198088
rect 54 197408 275435 197536
rect 880 196856 275435 197408
rect 54 196728 275435 196856
rect 880 196448 275435 196728
rect 54 196320 275435 196448
rect 880 195768 275435 196320
rect 54 195640 275435 195768
rect 880 195360 275435 195640
rect 54 195232 275435 195360
rect 880 194680 275435 195232
rect 54 194552 275435 194680
rect 880 194000 275435 194552
rect 54 193872 275435 194000
rect 880 193592 275435 193872
rect 54 193464 275435 193592
rect 880 192912 275435 193464
rect 54 192784 275435 192912
rect 880 192504 275435 192784
rect 54 192376 275435 192504
rect 880 191824 275435 192376
rect 54 191696 275435 191824
rect 880 191144 275435 191696
rect 54 191016 275435 191144
rect 880 190736 275435 191016
rect 54 190608 275435 190736
rect 880 190056 275435 190608
rect 54 189928 275435 190056
rect 880 189648 275435 189928
rect 54 189520 275435 189648
rect 880 188968 275435 189520
rect 54 188840 275435 188968
rect 880 188288 275435 188840
rect 54 188160 275435 188288
rect 880 187880 275435 188160
rect 54 187752 275435 187880
rect 880 187200 275435 187752
rect 54 187072 275435 187200
rect 880 186792 275435 187072
rect 54 186664 275435 186792
rect 880 186112 275435 186664
rect 54 185984 275435 186112
rect 880 185704 275435 185984
rect 54 185576 275435 185704
rect 880 185024 275435 185576
rect 54 184896 275435 185024
rect 880 184344 275435 184896
rect 54 184216 275435 184344
rect 880 183936 275435 184216
rect 54 183808 275435 183936
rect 880 183256 275435 183808
rect 54 183128 275435 183256
rect 880 182848 275435 183128
rect 54 182720 275435 182848
rect 880 182168 275435 182720
rect 54 182040 275435 182168
rect 880 181488 275435 182040
rect 54 181360 275435 181488
rect 880 181080 275435 181360
rect 54 180952 275435 181080
rect 880 180400 275435 180952
rect 54 180272 275435 180400
rect 880 179992 275435 180272
rect 54 179864 275435 179992
rect 880 179312 275435 179864
rect 54 179184 275435 179312
rect 880 178632 275435 179184
rect 54 178504 275435 178632
rect 880 178224 275435 178504
rect 54 178096 275435 178224
rect 880 177544 275435 178096
rect 54 177416 275435 177544
rect 880 177136 275435 177416
rect 54 177008 275435 177136
rect 880 176456 275435 177008
rect 54 176328 275435 176456
rect 880 175776 275435 176328
rect 54 175648 275435 175776
rect 880 175368 275435 175648
rect 54 175240 275435 175368
rect 880 174688 275435 175240
rect 54 174560 275435 174688
rect 880 174280 275435 174560
rect 54 174152 275435 174280
rect 880 173600 275435 174152
rect 54 173472 275435 173600
rect 880 172920 275435 173472
rect 54 172792 275435 172920
rect 880 172512 275435 172792
rect 54 172384 275435 172512
rect 880 171832 275435 172384
rect 54 171704 275435 171832
rect 880 171424 275435 171704
rect 54 171296 275435 171424
rect 880 170744 275435 171296
rect 54 170616 275435 170744
rect 880 170064 275435 170616
rect 54 169936 275435 170064
rect 880 169656 275435 169936
rect 54 169528 275435 169656
rect 880 168976 275435 169528
rect 54 168848 275435 168976
rect 880 168568 275435 168848
rect 54 168440 275435 168568
rect 880 167888 275435 168440
rect 54 167760 275435 167888
rect 880 167208 275435 167760
rect 54 167080 275435 167208
rect 880 166800 275435 167080
rect 54 166672 275435 166800
rect 880 166120 275435 166672
rect 54 165992 275435 166120
rect 880 165712 275435 165992
rect 54 165584 275435 165712
rect 880 165032 275435 165584
rect 54 164904 275435 165032
rect 880 164352 275435 164904
rect 54 164224 275435 164352
rect 880 163944 275435 164224
rect 54 163816 275435 163944
rect 880 163264 275435 163816
rect 54 163136 275435 163264
rect 880 162856 275435 163136
rect 54 162728 275435 162856
rect 880 162176 275435 162728
rect 54 162048 275435 162176
rect 880 161496 275435 162048
rect 54 161368 275435 161496
rect 880 161088 275435 161368
rect 54 160960 275435 161088
rect 880 160408 275435 160960
rect 54 160280 275435 160408
rect 880 160000 275435 160280
rect 54 159872 275435 160000
rect 880 159320 275435 159872
rect 54 159192 275435 159320
rect 880 158640 275435 159192
rect 54 158512 275435 158640
rect 880 158232 275435 158512
rect 54 158104 275435 158232
rect 880 157552 275435 158104
rect 54 157424 275435 157552
rect 880 157144 275435 157424
rect 54 157016 275435 157144
rect 880 156464 275435 157016
rect 54 156336 275435 156464
rect 880 155784 275435 156336
rect 54 155656 275435 155784
rect 880 155376 275435 155656
rect 54 155248 275435 155376
rect 880 154696 275435 155248
rect 54 154568 275435 154696
rect 880 154288 275435 154568
rect 54 154160 275435 154288
rect 880 153608 275435 154160
rect 54 153480 275435 153608
rect 880 152928 275435 153480
rect 54 152800 275435 152928
rect 880 152520 275435 152800
rect 54 152392 275435 152520
rect 880 151840 275435 152392
rect 54 151712 275435 151840
rect 880 151432 275435 151712
rect 54 151304 275435 151432
rect 880 150752 275435 151304
rect 54 150624 275435 150752
rect 880 150072 275435 150624
rect 54 149944 275435 150072
rect 880 149664 275435 149944
rect 54 149536 275435 149664
rect 880 148984 275435 149536
rect 54 148856 275435 148984
rect 880 148576 275435 148856
rect 54 148448 275435 148576
rect 880 147896 275435 148448
rect 54 147768 275435 147896
rect 880 147488 275435 147768
rect 54 147360 275435 147488
rect 880 146808 275435 147360
rect 54 146680 275435 146808
rect 880 146128 275435 146680
rect 54 146000 275435 146128
rect 880 145720 275435 146000
rect 54 145592 275435 145720
rect 880 145040 275435 145592
rect 54 144912 275435 145040
rect 880 144632 275435 144912
rect 54 144504 275435 144632
rect 880 143952 275435 144504
rect 54 143824 275435 143952
rect 880 143272 275435 143824
rect 54 143144 275435 143272
rect 880 142864 275435 143144
rect 54 142736 275435 142864
rect 880 142184 275435 142736
rect 54 142056 275435 142184
rect 880 141776 275435 142056
rect 54 141648 275435 141776
rect 880 141096 275435 141648
rect 54 140968 275435 141096
rect 880 140416 275435 140968
rect 54 140288 275435 140416
rect 880 140008 275435 140288
rect 54 139880 275435 140008
rect 880 139328 275435 139880
rect 54 139200 275435 139328
rect 880 138920 275435 139200
rect 54 138792 275435 138920
rect 880 138240 275435 138792
rect 54 138112 275435 138240
rect 880 137560 275435 138112
rect 54 137432 275435 137560
rect 880 137152 275435 137432
rect 54 137024 275435 137152
rect 880 136472 275435 137024
rect 54 136344 275435 136472
rect 880 136064 275435 136344
rect 54 135936 275435 136064
rect 880 135384 275435 135936
rect 54 135256 275435 135384
rect 880 134704 275435 135256
rect 54 134576 275435 134704
rect 880 134296 275435 134576
rect 54 134168 275435 134296
rect 880 133616 275435 134168
rect 54 133488 275435 133616
rect 880 133208 275435 133488
rect 54 133080 275435 133208
rect 880 132528 275435 133080
rect 54 132400 275435 132528
rect 880 131848 275435 132400
rect 54 131720 275435 131848
rect 880 131440 275435 131720
rect 54 131312 275435 131440
rect 880 130760 275435 131312
rect 54 130632 275435 130760
rect 880 130352 275435 130632
rect 54 130224 275435 130352
rect 880 129672 275435 130224
rect 54 129544 275435 129672
rect 880 128992 275435 129544
rect 54 128864 275435 128992
rect 880 128584 275435 128864
rect 54 128456 275435 128584
rect 880 127904 275435 128456
rect 54 127776 275435 127904
rect 880 127496 275435 127776
rect 54 127368 275435 127496
rect 880 126816 275435 127368
rect 54 126688 275435 126816
rect 880 126136 275435 126688
rect 54 126008 275435 126136
rect 880 125728 275435 126008
rect 54 125600 275435 125728
rect 880 125048 275435 125600
rect 54 124920 275435 125048
rect 880 124640 275435 124920
rect 54 124512 275435 124640
rect 880 123960 275435 124512
rect 54 123832 275435 123960
rect 880 123280 275435 123832
rect 54 123152 275435 123280
rect 880 122872 275435 123152
rect 54 122744 275435 122872
rect 880 122192 275435 122744
rect 54 122064 275435 122192
rect 880 121784 275435 122064
rect 54 121656 275435 121784
rect 880 121104 275435 121656
rect 54 120976 275435 121104
rect 880 120424 275435 120976
rect 54 120296 275435 120424
rect 880 120016 275435 120296
rect 54 119888 275435 120016
rect 880 119336 275435 119888
rect 54 119208 275435 119336
rect 880 118928 275435 119208
rect 54 118800 275435 118928
rect 880 118248 275435 118800
rect 54 118120 275435 118248
rect 880 117568 275435 118120
rect 54 117440 275435 117568
rect 880 117160 275435 117440
rect 54 117032 275435 117160
rect 880 116480 275435 117032
rect 54 116352 275435 116480
rect 880 116072 275435 116352
rect 54 115944 275435 116072
rect 880 115392 275435 115944
rect 54 115264 275435 115392
rect 880 114712 275435 115264
rect 54 114584 275435 114712
rect 880 114304 275435 114584
rect 54 114176 275435 114304
rect 880 113624 275435 114176
rect 54 113496 275435 113624
rect 880 113216 275435 113496
rect 54 113088 275435 113216
rect 880 112536 275435 113088
rect 54 112408 275435 112536
rect 880 112128 275435 112408
rect 54 112000 275435 112128
rect 880 111448 275435 112000
rect 54 111320 275435 111448
rect 880 110768 275435 111320
rect 54 110640 275435 110768
rect 880 110360 275435 110640
rect 54 110232 275435 110360
rect 880 109680 275435 110232
rect 54 109552 275435 109680
rect 880 109272 275435 109552
rect 54 109144 275435 109272
rect 880 108592 275435 109144
rect 54 108464 275435 108592
rect 880 107912 275435 108464
rect 54 107784 275435 107912
rect 880 107504 275435 107784
rect 54 107376 275435 107504
rect 880 106824 275435 107376
rect 54 106696 275435 106824
rect 880 106416 275435 106696
rect 54 106288 275435 106416
rect 880 105736 275435 106288
rect 54 105608 275435 105736
rect 880 105056 275435 105608
rect 54 104928 275435 105056
rect 880 104648 275435 104928
rect 54 104520 275435 104648
rect 880 103968 275435 104520
rect 54 103840 275435 103968
rect 880 103560 275435 103840
rect 54 103432 275435 103560
rect 880 102880 275435 103432
rect 54 102752 275435 102880
rect 880 102200 275435 102752
rect 54 102072 275435 102200
rect 880 101792 275435 102072
rect 54 101664 275435 101792
rect 880 101112 275435 101664
rect 54 100984 275435 101112
rect 880 100704 275435 100984
rect 54 100576 275435 100704
rect 880 100024 275435 100576
rect 54 99896 275435 100024
rect 880 99344 275435 99896
rect 54 99216 275435 99344
rect 880 98936 275435 99216
rect 54 98808 275435 98936
rect 880 98256 275435 98808
rect 54 98128 275435 98256
rect 880 97848 275435 98128
rect 54 97720 275435 97848
rect 880 97168 275435 97720
rect 54 97040 275435 97168
rect 880 96488 275435 97040
rect 54 96360 275435 96488
rect 880 96080 275435 96360
rect 54 95952 275435 96080
rect 880 95400 275435 95952
rect 54 95272 275435 95400
rect 880 94992 275435 95272
rect 54 94864 275435 94992
rect 880 94312 275435 94864
rect 54 94184 275435 94312
rect 880 93632 275435 94184
rect 54 93504 275435 93632
rect 880 93224 275435 93504
rect 54 93096 275435 93224
rect 880 92544 275435 93096
rect 54 92416 275435 92544
rect 880 92136 275435 92416
rect 54 92008 275435 92136
rect 880 91456 275435 92008
rect 54 91328 275435 91456
rect 880 90776 275435 91328
rect 54 90648 275435 90776
rect 880 90368 275435 90648
rect 54 90240 275435 90368
rect 880 89688 275435 90240
rect 54 89560 275435 89688
rect 880 89280 275435 89560
rect 54 89152 275435 89280
rect 880 88600 275435 89152
rect 54 88472 275435 88600
rect 880 87920 275435 88472
rect 54 87792 275435 87920
rect 880 87512 275435 87792
rect 54 87384 275435 87512
rect 880 86832 275435 87384
rect 54 86704 275435 86832
rect 880 86424 275435 86704
rect 54 86296 275435 86424
rect 880 85744 275435 86296
rect 54 85616 275435 85744
rect 880 85064 275435 85616
rect 54 84936 275435 85064
rect 880 84656 275435 84936
rect 54 84528 275435 84656
rect 880 83976 275435 84528
rect 54 83848 275435 83976
rect 880 83568 275435 83848
rect 54 83440 275435 83568
rect 880 82888 275435 83440
rect 54 82760 275435 82888
rect 880 82208 275435 82760
rect 54 82080 275435 82208
rect 880 81800 275435 82080
rect 54 81672 275435 81800
rect 880 81120 275435 81672
rect 54 80992 275435 81120
rect 880 80712 275435 80992
rect 54 80584 275435 80712
rect 880 80032 275435 80584
rect 54 79904 275435 80032
rect 880 79352 275435 79904
rect 54 79224 275435 79352
rect 880 78944 275435 79224
rect 54 78816 275435 78944
rect 880 78264 275435 78816
rect 54 78136 275435 78264
rect 880 77856 275435 78136
rect 54 77728 275435 77856
rect 880 77176 275435 77728
rect 54 77048 275435 77176
rect 880 76496 275435 77048
rect 54 76368 275435 76496
rect 880 76088 275435 76368
rect 54 75960 275435 76088
rect 880 75408 275435 75960
rect 54 75280 275435 75408
rect 880 75000 275435 75280
rect 54 74872 275435 75000
rect 880 74320 275435 74872
rect 54 74192 275435 74320
rect 880 73912 275435 74192
rect 54 73784 275435 73912
rect 880 73232 275435 73784
rect 54 73104 275435 73232
rect 880 72552 275435 73104
rect 54 72424 275435 72552
rect 880 72144 275435 72424
rect 54 72016 275435 72144
rect 880 71464 275435 72016
rect 54 71336 275435 71464
rect 880 71056 275435 71336
rect 54 70928 275435 71056
rect 880 70376 275435 70928
rect 54 70248 275435 70376
rect 880 69696 275435 70248
rect 54 69568 275435 69696
rect 880 69288 275435 69568
rect 54 69160 275435 69288
rect 880 68608 275435 69160
rect 54 68480 275435 68608
rect 880 68200 275435 68480
rect 54 68072 275435 68200
rect 880 67520 275435 68072
rect 54 67392 275435 67520
rect 880 66840 275435 67392
rect 54 66712 275435 66840
rect 880 66432 275435 66712
rect 54 66304 275435 66432
rect 880 65752 275435 66304
rect 54 65624 275435 65752
rect 880 65344 275435 65624
rect 54 65216 275435 65344
rect 880 64664 275435 65216
rect 54 64536 275435 64664
rect 880 63984 275435 64536
rect 54 63856 275435 63984
rect 880 63576 275435 63856
rect 54 63448 275435 63576
rect 880 62896 275435 63448
rect 54 62768 275435 62896
rect 880 62488 275435 62768
rect 54 62360 275435 62488
rect 880 61808 275435 62360
rect 54 61680 275435 61808
rect 880 61128 275435 61680
rect 54 61000 275435 61128
rect 880 60720 275435 61000
rect 54 60592 275435 60720
rect 880 60040 275435 60592
rect 54 59912 275435 60040
rect 880 59632 275435 59912
rect 54 59504 275435 59632
rect 880 58952 275435 59504
rect 54 58824 275435 58952
rect 880 58272 275435 58824
rect 54 58144 275435 58272
rect 880 57864 275435 58144
rect 54 57736 275435 57864
rect 880 57184 275435 57736
rect 54 57056 275435 57184
rect 880 56776 275435 57056
rect 54 56648 275435 56776
rect 880 56096 275435 56648
rect 54 55968 275435 56096
rect 880 55416 275435 55968
rect 54 55288 275435 55416
rect 880 55008 275435 55288
rect 54 54880 275435 55008
rect 880 54328 275435 54880
rect 54 54200 275435 54328
rect 880 53920 275435 54200
rect 54 53792 275435 53920
rect 880 53240 275435 53792
rect 54 53112 275435 53240
rect 880 52560 275435 53112
rect 54 52432 275435 52560
rect 880 52152 275435 52432
rect 54 52024 275435 52152
rect 880 51472 275435 52024
rect 54 51344 275435 51472
rect 880 51064 275435 51344
rect 54 50936 275435 51064
rect 880 50384 275435 50936
rect 54 50256 275435 50384
rect 880 49704 275435 50256
rect 54 49576 275435 49704
rect 880 49296 275435 49576
rect 54 49168 275435 49296
rect 880 48616 275435 49168
rect 54 48488 275435 48616
rect 880 48208 275435 48488
rect 54 48080 275435 48208
rect 880 47528 275435 48080
rect 54 47400 275435 47528
rect 880 46848 275435 47400
rect 54 46720 275435 46848
rect 880 46440 275435 46720
rect 54 46312 275435 46440
rect 880 45760 275435 46312
rect 54 45632 275435 45760
rect 880 45352 275435 45632
rect 54 45224 275435 45352
rect 880 44672 275435 45224
rect 54 44544 275435 44672
rect 880 43992 275435 44544
rect 54 43864 275435 43992
rect 880 43584 275435 43864
rect 54 43456 275435 43584
rect 880 42904 275435 43456
rect 54 42776 275435 42904
rect 880 42496 275435 42776
rect 54 42368 275435 42496
rect 880 41816 275435 42368
rect 54 41688 275435 41816
rect 880 41136 275435 41688
rect 54 41008 275435 41136
rect 880 40728 275435 41008
rect 54 40600 275435 40728
rect 880 40048 275435 40600
rect 54 39920 275435 40048
rect 880 39640 275435 39920
rect 54 39512 275435 39640
rect 880 38960 275435 39512
rect 54 38832 275435 38960
rect 880 38280 275435 38832
rect 54 38152 275435 38280
rect 880 37872 275435 38152
rect 54 37744 275435 37872
rect 880 37192 275435 37744
rect 54 37064 275435 37192
rect 880 36784 275435 37064
rect 54 36656 275435 36784
rect 880 36104 275435 36656
rect 54 35976 275435 36104
rect 880 35696 275435 35976
rect 54 35568 275435 35696
rect 880 35016 275435 35568
rect 54 34888 275435 35016
rect 880 34336 275435 34888
rect 54 34208 275435 34336
rect 880 33928 275435 34208
rect 54 33800 275435 33928
rect 880 33248 275435 33800
rect 54 33120 275435 33248
rect 880 32840 275435 33120
rect 54 32712 275435 32840
rect 880 32160 275435 32712
rect 54 32032 275435 32160
rect 880 31480 275435 32032
rect 54 31352 275435 31480
rect 880 31072 275435 31352
rect 54 30944 275435 31072
rect 880 30392 275435 30944
rect 54 30264 275435 30392
rect 880 29984 275435 30264
rect 54 29856 275435 29984
rect 880 29304 275435 29856
rect 54 29176 275435 29304
rect 880 28624 275435 29176
rect 54 28496 275435 28624
rect 880 28216 275435 28496
rect 54 28088 275435 28216
rect 880 27536 275435 28088
rect 54 27408 275435 27536
rect 880 27128 275435 27408
rect 54 27000 275435 27128
rect 880 26448 275435 27000
rect 54 26320 275435 26448
rect 880 25768 275435 26320
rect 54 25640 275435 25768
rect 880 25360 275435 25640
rect 54 25232 275435 25360
rect 880 24680 275435 25232
rect 54 24552 275435 24680
rect 880 24272 275435 24552
rect 54 24144 275435 24272
rect 880 23592 275435 24144
rect 54 23464 275435 23592
rect 880 22912 275435 23464
rect 54 22784 275435 22912
rect 880 22504 275435 22784
rect 54 22376 275435 22504
rect 880 21824 275435 22376
rect 54 21696 275435 21824
rect 880 21416 275435 21696
rect 54 21288 275435 21416
rect 880 20736 275435 21288
rect 54 20608 275435 20736
rect 880 20056 275435 20608
rect 54 19928 275435 20056
rect 880 19648 275435 19928
rect 54 19520 275435 19648
rect 880 18968 275435 19520
rect 54 18840 275435 18968
rect 880 18560 275435 18840
rect 54 18432 275435 18560
rect 880 17880 275435 18432
rect 54 17752 275435 17880
rect 880 17200 275435 17752
rect 54 17072 275435 17200
rect 880 16792 275435 17072
rect 54 16664 275435 16792
rect 880 16112 275435 16664
rect 54 15984 275435 16112
rect 880 15704 275435 15984
rect 54 15576 275435 15704
rect 880 15024 275435 15576
rect 54 14896 275435 15024
rect 880 14344 275435 14896
rect 54 14216 275435 14344
rect 880 13936 275435 14216
rect 54 13808 275435 13936
rect 880 13256 275435 13808
rect 54 13128 275435 13256
rect 880 12848 275435 13128
rect 54 12720 275435 12848
rect 880 12168 275435 12720
rect 54 12040 275435 12168
rect 880 11488 275435 12040
rect 54 11360 275435 11488
rect 880 11080 275435 11360
rect 54 10952 275435 11080
rect 880 10400 275435 10952
rect 54 10272 275435 10400
rect 880 9992 275435 10272
rect 54 9864 275435 9992
rect 880 9312 275435 9864
rect 54 9184 275435 9312
rect 880 8632 275435 9184
rect 54 8504 275435 8632
rect 880 8224 275435 8504
rect 54 8096 275435 8224
rect 880 7544 275435 8096
rect 54 7416 275435 7544
rect 880 7136 275435 7416
rect 54 7008 275435 7136
rect 880 6456 275435 7008
rect 54 6328 275435 6456
rect 880 5776 275435 6328
rect 54 5648 275435 5776
rect 880 5368 275435 5648
rect 54 5240 275435 5368
rect 880 4688 275435 5240
rect 54 4560 275435 4688
rect 880 4280 275435 4560
rect 54 4152 275435 4280
rect 880 3600 275435 4152
rect 54 3472 275435 3600
rect 880 2920 275435 3472
rect 54 2792 275435 2920
rect 880 2512 275435 2792
rect 54 2384 275435 2512
rect 880 1832 275435 2384
rect 54 1704 275435 1832
rect 880 1424 275435 1704
rect 54 1296 275435 1424
rect 880 744 275435 1296
rect 54 616 275435 744
rect 880 171 275435 616
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
rect 111728 2128 112048 297616
rect 127088 2128 127408 297616
rect 142448 2128 142768 297616
rect 157808 2128 158128 297616
rect 173168 2128 173488 297616
rect 188528 2128 188848 297616
rect 203888 2128 204208 297616
rect 219248 2128 219568 297616
rect 234608 2128 234928 297616
rect 249968 2128 250288 297616
rect 265328 2128 265648 297616
<< obsm4 >>
rect 59 297696 273549 299437
rect 59 2048 4128 297696
rect 4608 2048 19488 297696
rect 19968 2048 34848 297696
rect 35328 2048 50208 297696
rect 50688 2048 65568 297696
rect 66048 2048 80928 297696
rect 81408 2048 96288 297696
rect 96768 2048 111648 297696
rect 112128 2048 127008 297696
rect 127488 2048 142368 297696
rect 142848 2048 157728 297696
rect 158208 2048 173088 297696
rect 173568 2048 188448 297696
rect 188928 2048 203808 297696
rect 204288 2048 219168 297696
rect 219648 2048 234528 297696
rect 235008 2048 249888 297696
rect 250368 2048 265248 297696
rect 265728 2048 273549 297696
rect 59 1803 273549 2048
<< labels >>
rlabel metal2 s 478 0 534 800 6 clk
port 1 nsew signal input
rlabel metal3 s 0 247936 800 248056 6 core_id[0]
port 2 nsew signal input
rlabel metal3 s 0 251472 800 251592 6 core_id[10]
port 3 nsew signal input
rlabel metal3 s 0 251880 800 252000 6 core_id[11]
port 4 nsew signal input
rlabel metal3 s 0 252288 800 252408 6 core_id[12]
port 5 nsew signal input
rlabel metal3 s 0 252560 800 252680 6 core_id[13]
port 6 nsew signal input
rlabel metal3 s 0 252968 800 253088 6 core_id[14]
port 7 nsew signal input
rlabel metal3 s 0 253240 800 253360 6 core_id[15]
port 8 nsew signal input
rlabel metal3 s 0 253648 800 253768 6 core_id[16]
port 9 nsew signal input
rlabel metal3 s 0 254056 800 254176 6 core_id[17]
port 10 nsew signal input
rlabel metal3 s 0 254328 800 254448 6 core_id[18]
port 11 nsew signal input
rlabel metal3 s 0 254736 800 254856 6 core_id[19]
port 12 nsew signal input
rlabel metal3 s 0 248344 800 248464 6 core_id[1]
port 13 nsew signal input
rlabel metal3 s 0 255144 800 255264 6 core_id[20]
port 14 nsew signal input
rlabel metal3 s 0 255416 800 255536 6 core_id[21]
port 15 nsew signal input
rlabel metal3 s 0 255824 800 255944 6 core_id[22]
port 16 nsew signal input
rlabel metal3 s 0 256096 800 256216 6 core_id[23]
port 17 nsew signal input
rlabel metal3 s 0 256504 800 256624 6 core_id[24]
port 18 nsew signal input
rlabel metal3 s 0 256912 800 257032 6 core_id[25]
port 19 nsew signal input
rlabel metal3 s 0 257184 800 257304 6 core_id[26]
port 20 nsew signal input
rlabel metal3 s 0 257592 800 257712 6 core_id[27]
port 21 nsew signal input
rlabel metal3 s 0 248616 800 248736 6 core_id[2]
port 22 nsew signal input
rlabel metal3 s 0 249024 800 249144 6 core_id[3]
port 23 nsew signal input
rlabel metal3 s 0 249432 800 249552 6 core_id[4]
port 24 nsew signal input
rlabel metal3 s 0 249704 800 249824 6 core_id[5]
port 25 nsew signal input
rlabel metal3 s 0 250112 800 250232 6 core_id[6]
port 26 nsew signal input
rlabel metal3 s 0 250384 800 250504 6 core_id[7]
port 27 nsew signal input
rlabel metal3 s 0 250792 800 250912 6 core_id[8]
port 28 nsew signal input
rlabel metal3 s 0 251200 800 251320 6 core_id[9]
port 29 nsew signal input
rlabel metal3 s 0 173000 800 173120 6 dbg_bus_clk_en
port 30 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 dbg_rst_l
port 31 nsew signal input
rlabel metal3 s 0 173680 800 173800 6 dccm_ext_in_pkt[0]
port 32 nsew signal input
rlabel metal3 s 0 177216 800 177336 6 dccm_ext_in_pkt[10]
port 33 nsew signal input
rlabel metal3 s 0 177624 800 177744 6 dccm_ext_in_pkt[11]
port 34 nsew signal input
rlabel metal3 s 0 177896 800 178016 6 dccm_ext_in_pkt[12]
port 35 nsew signal input
rlabel metal3 s 0 178304 800 178424 6 dccm_ext_in_pkt[13]
port 36 nsew signal input
rlabel metal3 s 0 178712 800 178832 6 dccm_ext_in_pkt[14]
port 37 nsew signal input
rlabel metal3 s 0 178984 800 179104 6 dccm_ext_in_pkt[15]
port 38 nsew signal input
rlabel metal3 s 0 179392 800 179512 6 dccm_ext_in_pkt[16]
port 39 nsew signal input
rlabel metal3 s 0 179664 800 179784 6 dccm_ext_in_pkt[17]
port 40 nsew signal input
rlabel metal3 s 0 180072 800 180192 6 dccm_ext_in_pkt[18]
port 41 nsew signal input
rlabel metal3 s 0 180480 800 180600 6 dccm_ext_in_pkt[19]
port 42 nsew signal input
rlabel metal3 s 0 173952 800 174072 6 dccm_ext_in_pkt[1]
port 43 nsew signal input
rlabel metal3 s 0 180752 800 180872 6 dccm_ext_in_pkt[20]
port 44 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 dccm_ext_in_pkt[21]
port 45 nsew signal input
rlabel metal3 s 0 181568 800 181688 6 dccm_ext_in_pkt[22]
port 46 nsew signal input
rlabel metal3 s 0 181840 800 181960 6 dccm_ext_in_pkt[23]
port 47 nsew signal input
rlabel metal3 s 0 182248 800 182368 6 dccm_ext_in_pkt[24]
port 48 nsew signal input
rlabel metal3 s 0 182520 800 182640 6 dccm_ext_in_pkt[25]
port 49 nsew signal input
rlabel metal3 s 0 182928 800 183048 6 dccm_ext_in_pkt[26]
port 50 nsew signal input
rlabel metal3 s 0 183336 800 183456 6 dccm_ext_in_pkt[27]
port 51 nsew signal input
rlabel metal3 s 0 183608 800 183728 6 dccm_ext_in_pkt[28]
port 52 nsew signal input
rlabel metal3 s 0 184016 800 184136 6 dccm_ext_in_pkt[29]
port 53 nsew signal input
rlabel metal3 s 0 174360 800 174480 6 dccm_ext_in_pkt[2]
port 54 nsew signal input
rlabel metal3 s 0 184424 800 184544 6 dccm_ext_in_pkt[30]
port 55 nsew signal input
rlabel metal3 s 0 184696 800 184816 6 dccm_ext_in_pkt[31]
port 56 nsew signal input
rlabel metal3 s 0 185104 800 185224 6 dccm_ext_in_pkt[32]
port 57 nsew signal input
rlabel metal3 s 0 185376 800 185496 6 dccm_ext_in_pkt[33]
port 58 nsew signal input
rlabel metal3 s 0 185784 800 185904 6 dccm_ext_in_pkt[34]
port 59 nsew signal input
rlabel metal3 s 0 186192 800 186312 6 dccm_ext_in_pkt[35]
port 60 nsew signal input
rlabel metal3 s 0 186464 800 186584 6 dccm_ext_in_pkt[36]
port 61 nsew signal input
rlabel metal3 s 0 186872 800 186992 6 dccm_ext_in_pkt[37]
port 62 nsew signal input
rlabel metal3 s 0 187280 800 187400 6 dccm_ext_in_pkt[38]
port 63 nsew signal input
rlabel metal3 s 0 187552 800 187672 6 dccm_ext_in_pkt[39]
port 64 nsew signal input
rlabel metal3 s 0 174768 800 174888 6 dccm_ext_in_pkt[3]
port 65 nsew signal input
rlabel metal3 s 0 187960 800 188080 6 dccm_ext_in_pkt[40]
port 66 nsew signal input
rlabel metal3 s 0 188368 800 188488 6 dccm_ext_in_pkt[41]
port 67 nsew signal input
rlabel metal3 s 0 188640 800 188760 6 dccm_ext_in_pkt[42]
port 68 nsew signal input
rlabel metal3 s 0 189048 800 189168 6 dccm_ext_in_pkt[43]
port 69 nsew signal input
rlabel metal3 s 0 189320 800 189440 6 dccm_ext_in_pkt[44]
port 70 nsew signal input
rlabel metal3 s 0 189728 800 189848 6 dccm_ext_in_pkt[45]
port 71 nsew signal input
rlabel metal3 s 0 190136 800 190256 6 dccm_ext_in_pkt[46]
port 72 nsew signal input
rlabel metal3 s 0 190408 800 190528 6 dccm_ext_in_pkt[47]
port 73 nsew signal input
rlabel metal3 s 0 175040 800 175160 6 dccm_ext_in_pkt[4]
port 74 nsew signal input
rlabel metal3 s 0 175448 800 175568 6 dccm_ext_in_pkt[5]
port 75 nsew signal input
rlabel metal3 s 0 175856 800 175976 6 dccm_ext_in_pkt[6]
port 76 nsew signal input
rlabel metal3 s 0 176128 800 176248 6 dccm_ext_in_pkt[7]
port 77 nsew signal input
rlabel metal3 s 0 176536 800 176656 6 dccm_ext_in_pkt[8]
port 78 nsew signal input
rlabel metal3 s 0 176808 800 176928 6 dccm_ext_in_pkt[9]
port 79 nsew signal input
rlabel metal3 s 0 259768 800 259888 6 debug_brkpt_status
port 80 nsew signal output
rlabel metal3 s 0 233656 800 233776 6 dec_tlu_perfcnt0
port 81 nsew signal output
rlabel metal3 s 0 234064 800 234184 6 dec_tlu_perfcnt1
port 82 nsew signal output
rlabel metal3 s 0 234336 800 234456 6 dec_tlu_perfcnt2
port 83 nsew signal output
rlabel metal3 s 0 234744 800 234864 6 dec_tlu_perfcnt3
port 84 nsew signal output
rlabel metal3 s 0 173272 800 173392 6 dma_bus_clk_en
port 85 nsew signal input
rlabel metal3 s 0 108944 800 109064 6 dma_haddr[0]
port 86 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 dma_haddr[10]
port 87 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 dma_haddr[11]
port 88 nsew signal input
rlabel metal3 s 0 113296 800 113416 6 dma_haddr[12]
port 89 nsew signal input
rlabel metal3 s 0 113704 800 113824 6 dma_haddr[13]
port 90 nsew signal input
rlabel metal3 s 0 113976 800 114096 6 dma_haddr[14]
port 91 nsew signal input
rlabel metal3 s 0 114384 800 114504 6 dma_haddr[15]
port 92 nsew signal input
rlabel metal3 s 0 114792 800 114912 6 dma_haddr[16]
port 93 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 dma_haddr[17]
port 94 nsew signal input
rlabel metal3 s 0 115472 800 115592 6 dma_haddr[18]
port 95 nsew signal input
rlabel metal3 s 0 115744 800 115864 6 dma_haddr[19]
port 96 nsew signal input
rlabel metal3 s 0 109352 800 109472 6 dma_haddr[1]
port 97 nsew signal input
rlabel metal3 s 0 116152 800 116272 6 dma_haddr[20]
port 98 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 dma_haddr[21]
port 99 nsew signal input
rlabel metal3 s 0 116832 800 116952 6 dma_haddr[22]
port 100 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 dma_haddr[23]
port 101 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 dma_haddr[24]
port 102 nsew signal input
rlabel metal3 s 0 117920 800 118040 6 dma_haddr[25]
port 103 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 dma_haddr[26]
port 104 nsew signal input
rlabel metal3 s 0 118600 800 118720 6 dma_haddr[27]
port 105 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 dma_haddr[28]
port 106 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 dma_haddr[29]
port 107 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 dma_haddr[2]
port 108 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 dma_haddr[30]
port 109 nsew signal input
rlabel metal3 s 0 120096 800 120216 6 dma_haddr[31]
port 110 nsew signal input
rlabel metal3 s 0 110032 800 110152 6 dma_haddr[3]
port 111 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 dma_haddr[4]
port 112 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 dma_haddr[5]
port 113 nsew signal input
rlabel metal3 s 0 111120 800 111240 6 dma_haddr[6]
port 114 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 dma_haddr[7]
port 115 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 dma_haddr[8]
port 116 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 dma_haddr[9]
port 117 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 dma_hburst[0]
port 118 nsew signal input
rlabel metal3 s 0 120776 800 120896 6 dma_hburst[1]
port 119 nsew signal input
rlabel metal3 s 0 121184 800 121304 6 dma_hburst[2]
port 120 nsew signal input
rlabel metal3 s 0 121456 800 121576 6 dma_hmastlock
port 121 nsew signal input
rlabel metal3 s 0 121864 800 121984 6 dma_hprot[0]
port 122 nsew signal input
rlabel metal3 s 0 122272 800 122392 6 dma_hprot[1]
port 123 nsew signal input
rlabel metal3 s 0 122544 800 122664 6 dma_hprot[2]
port 124 nsew signal input
rlabel metal3 s 0 122952 800 123072 6 dma_hprot[3]
port 125 nsew signal input
rlabel metal3 s 0 148656 800 148776 6 dma_hrdata[0]
port 126 nsew signal output
rlabel metal3 s 0 152192 800 152312 6 dma_hrdata[10]
port 127 nsew signal output
rlabel metal3 s 0 152600 800 152720 6 dma_hrdata[11]
port 128 nsew signal output
rlabel metal3 s 0 153008 800 153128 6 dma_hrdata[12]
port 129 nsew signal output
rlabel metal3 s 0 153280 800 153400 6 dma_hrdata[13]
port 130 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 dma_hrdata[14]
port 131 nsew signal output
rlabel metal3 s 0 153960 800 154080 6 dma_hrdata[15]
port 132 nsew signal output
rlabel metal3 s 0 154368 800 154488 6 dma_hrdata[16]
port 133 nsew signal output
rlabel metal3 s 0 154776 800 154896 6 dma_hrdata[17]
port 134 nsew signal output
rlabel metal3 s 0 155048 800 155168 6 dma_hrdata[18]
port 135 nsew signal output
rlabel metal3 s 0 155456 800 155576 6 dma_hrdata[19]
port 136 nsew signal output
rlabel metal3 s 0 149064 800 149184 6 dma_hrdata[1]
port 137 nsew signal output
rlabel metal3 s 0 155864 800 155984 6 dma_hrdata[20]
port 138 nsew signal output
rlabel metal3 s 0 156136 800 156256 6 dma_hrdata[21]
port 139 nsew signal output
rlabel metal3 s 0 156544 800 156664 6 dma_hrdata[22]
port 140 nsew signal output
rlabel metal3 s 0 156816 800 156936 6 dma_hrdata[23]
port 141 nsew signal output
rlabel metal3 s 0 157224 800 157344 6 dma_hrdata[24]
port 142 nsew signal output
rlabel metal3 s 0 157632 800 157752 6 dma_hrdata[25]
port 143 nsew signal output
rlabel metal3 s 0 157904 800 158024 6 dma_hrdata[26]
port 144 nsew signal output
rlabel metal3 s 0 158312 800 158432 6 dma_hrdata[27]
port 145 nsew signal output
rlabel metal3 s 0 158720 800 158840 6 dma_hrdata[28]
port 146 nsew signal output
rlabel metal3 s 0 158992 800 159112 6 dma_hrdata[29]
port 147 nsew signal output
rlabel metal3 s 0 149336 800 149456 6 dma_hrdata[2]
port 148 nsew signal output
rlabel metal3 s 0 159400 800 159520 6 dma_hrdata[30]
port 149 nsew signal output
rlabel metal3 s 0 159672 800 159792 6 dma_hrdata[31]
port 150 nsew signal output
rlabel metal3 s 0 160080 800 160200 6 dma_hrdata[32]
port 151 nsew signal output
rlabel metal3 s 0 160488 800 160608 6 dma_hrdata[33]
port 152 nsew signal output
rlabel metal3 s 0 160760 800 160880 6 dma_hrdata[34]
port 153 nsew signal output
rlabel metal3 s 0 161168 800 161288 6 dma_hrdata[35]
port 154 nsew signal output
rlabel metal3 s 0 161576 800 161696 6 dma_hrdata[36]
port 155 nsew signal output
rlabel metal3 s 0 161848 800 161968 6 dma_hrdata[37]
port 156 nsew signal output
rlabel metal3 s 0 162256 800 162376 6 dma_hrdata[38]
port 157 nsew signal output
rlabel metal3 s 0 162528 800 162648 6 dma_hrdata[39]
port 158 nsew signal output
rlabel metal3 s 0 149744 800 149864 6 dma_hrdata[3]
port 159 nsew signal output
rlabel metal3 s 0 162936 800 163056 6 dma_hrdata[40]
port 160 nsew signal output
rlabel metal3 s 0 163344 800 163464 6 dma_hrdata[41]
port 161 nsew signal output
rlabel metal3 s 0 163616 800 163736 6 dma_hrdata[42]
port 162 nsew signal output
rlabel metal3 s 0 164024 800 164144 6 dma_hrdata[43]
port 163 nsew signal output
rlabel metal3 s 0 164432 800 164552 6 dma_hrdata[44]
port 164 nsew signal output
rlabel metal3 s 0 164704 800 164824 6 dma_hrdata[45]
port 165 nsew signal output
rlabel metal3 s 0 165112 800 165232 6 dma_hrdata[46]
port 166 nsew signal output
rlabel metal3 s 0 165384 800 165504 6 dma_hrdata[47]
port 167 nsew signal output
rlabel metal3 s 0 165792 800 165912 6 dma_hrdata[48]
port 168 nsew signal output
rlabel metal3 s 0 166200 800 166320 6 dma_hrdata[49]
port 169 nsew signal output
rlabel metal3 s 0 150152 800 150272 6 dma_hrdata[4]
port 170 nsew signal output
rlabel metal3 s 0 166472 800 166592 6 dma_hrdata[50]
port 171 nsew signal output
rlabel metal3 s 0 166880 800 167000 6 dma_hrdata[51]
port 172 nsew signal output
rlabel metal3 s 0 167288 800 167408 6 dma_hrdata[52]
port 173 nsew signal output
rlabel metal3 s 0 167560 800 167680 6 dma_hrdata[53]
port 174 nsew signal output
rlabel metal3 s 0 167968 800 168088 6 dma_hrdata[54]
port 175 nsew signal output
rlabel metal3 s 0 168240 800 168360 6 dma_hrdata[55]
port 176 nsew signal output
rlabel metal3 s 0 168648 800 168768 6 dma_hrdata[56]
port 177 nsew signal output
rlabel metal3 s 0 169056 800 169176 6 dma_hrdata[57]
port 178 nsew signal output
rlabel metal3 s 0 169328 800 169448 6 dma_hrdata[58]
port 179 nsew signal output
rlabel metal3 s 0 169736 800 169856 6 dma_hrdata[59]
port 180 nsew signal output
rlabel metal3 s 0 150424 800 150544 6 dma_hrdata[5]
port 181 nsew signal output
rlabel metal3 s 0 170144 800 170264 6 dma_hrdata[60]
port 182 nsew signal output
rlabel metal3 s 0 170416 800 170536 6 dma_hrdata[61]
port 183 nsew signal output
rlabel metal3 s 0 170824 800 170944 6 dma_hrdata[62]
port 184 nsew signal output
rlabel metal3 s 0 171096 800 171216 6 dma_hrdata[63]
port 185 nsew signal output
rlabel metal3 s 0 150832 800 150952 6 dma_hrdata[6]
port 186 nsew signal output
rlabel metal3 s 0 151104 800 151224 6 dma_hrdata[7]
port 187 nsew signal output
rlabel metal3 s 0 151512 800 151632 6 dma_hrdata[8]
port 188 nsew signal output
rlabel metal3 s 0 151920 800 152040 6 dma_hrdata[9]
port 189 nsew signal output
rlabel metal3 s 0 148248 800 148368 6 dma_hreadyin
port 190 nsew signal input
rlabel metal3 s 0 171504 800 171624 6 dma_hreadyout
port 191 nsew signal output
rlabel metal3 s 0 171912 800 172032 6 dma_hresp
port 192 nsew signal output
rlabel metal3 s 0 108672 800 108792 6 dma_hsel
port 193 nsew signal input
rlabel metal3 s 0 123360 800 123480 6 dma_hsize[0]
port 194 nsew signal input
rlabel metal3 s 0 123632 800 123752 6 dma_hsize[1]
port 195 nsew signal input
rlabel metal3 s 0 124040 800 124160 6 dma_hsize[2]
port 196 nsew signal input
rlabel metal3 s 0 124312 800 124432 6 dma_htrans[0]
port 197 nsew signal input
rlabel metal3 s 0 124720 800 124840 6 dma_htrans[1]
port 198 nsew signal input
rlabel metal3 s 0 125400 800 125520 6 dma_hwdata[0]
port 199 nsew signal input
rlabel metal3 s 0 129072 800 129192 6 dma_hwdata[10]
port 200 nsew signal input
rlabel metal3 s 0 129344 800 129464 6 dma_hwdata[11]
port 201 nsew signal input
rlabel metal3 s 0 129752 800 129872 6 dma_hwdata[12]
port 202 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 dma_hwdata[13]
port 203 nsew signal input
rlabel metal3 s 0 130432 800 130552 6 dma_hwdata[14]
port 204 nsew signal input
rlabel metal3 s 0 130840 800 130960 6 dma_hwdata[15]
port 205 nsew signal input
rlabel metal3 s 0 131112 800 131232 6 dma_hwdata[16]
port 206 nsew signal input
rlabel metal3 s 0 131520 800 131640 6 dma_hwdata[17]
port 207 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 dma_hwdata[18]
port 208 nsew signal input
rlabel metal3 s 0 132200 800 132320 6 dma_hwdata[19]
port 209 nsew signal input
rlabel metal3 s 0 125808 800 125928 6 dma_hwdata[1]
port 210 nsew signal input
rlabel metal3 s 0 132608 800 132728 6 dma_hwdata[20]
port 211 nsew signal input
rlabel metal3 s 0 132880 800 133000 6 dma_hwdata[21]
port 212 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 dma_hwdata[22]
port 213 nsew signal input
rlabel metal3 s 0 133696 800 133816 6 dma_hwdata[23]
port 214 nsew signal input
rlabel metal3 s 0 133968 800 134088 6 dma_hwdata[24]
port 215 nsew signal input
rlabel metal3 s 0 134376 800 134496 6 dma_hwdata[25]
port 216 nsew signal input
rlabel metal3 s 0 134784 800 134904 6 dma_hwdata[26]
port 217 nsew signal input
rlabel metal3 s 0 135056 800 135176 6 dma_hwdata[27]
port 218 nsew signal input
rlabel metal3 s 0 135464 800 135584 6 dma_hwdata[28]
port 219 nsew signal input
rlabel metal3 s 0 135736 800 135856 6 dma_hwdata[29]
port 220 nsew signal input
rlabel metal3 s 0 126216 800 126336 6 dma_hwdata[2]
port 221 nsew signal input
rlabel metal3 s 0 136144 800 136264 6 dma_hwdata[30]
port 222 nsew signal input
rlabel metal3 s 0 136552 800 136672 6 dma_hwdata[31]
port 223 nsew signal input
rlabel metal3 s 0 136824 800 136944 6 dma_hwdata[32]
port 224 nsew signal input
rlabel metal3 s 0 137232 800 137352 6 dma_hwdata[33]
port 225 nsew signal input
rlabel metal3 s 0 137640 800 137760 6 dma_hwdata[34]
port 226 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 dma_hwdata[35]
port 227 nsew signal input
rlabel metal3 s 0 138320 800 138440 6 dma_hwdata[36]
port 228 nsew signal input
rlabel metal3 s 0 138592 800 138712 6 dma_hwdata[37]
port 229 nsew signal input
rlabel metal3 s 0 139000 800 139120 6 dma_hwdata[38]
port 230 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 dma_hwdata[39]
port 231 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 dma_hwdata[3]
port 232 nsew signal input
rlabel metal3 s 0 139680 800 139800 6 dma_hwdata[40]
port 233 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 dma_hwdata[41]
port 234 nsew signal input
rlabel metal3 s 0 140496 800 140616 6 dma_hwdata[42]
port 235 nsew signal input
rlabel metal3 s 0 140768 800 140888 6 dma_hwdata[43]
port 236 nsew signal input
rlabel metal3 s 0 141176 800 141296 6 dma_hwdata[44]
port 237 nsew signal input
rlabel metal3 s 0 141448 800 141568 6 dma_hwdata[45]
port 238 nsew signal input
rlabel metal3 s 0 141856 800 141976 6 dma_hwdata[46]
port 239 nsew signal input
rlabel metal3 s 0 142264 800 142384 6 dma_hwdata[47]
port 240 nsew signal input
rlabel metal3 s 0 142536 800 142656 6 dma_hwdata[48]
port 241 nsew signal input
rlabel metal3 s 0 142944 800 143064 6 dma_hwdata[49]
port 242 nsew signal input
rlabel metal3 s 0 126896 800 127016 6 dma_hwdata[4]
port 243 nsew signal input
rlabel metal3 s 0 143352 800 143472 6 dma_hwdata[50]
port 244 nsew signal input
rlabel metal3 s 0 143624 800 143744 6 dma_hwdata[51]
port 245 nsew signal input
rlabel metal3 s 0 144032 800 144152 6 dma_hwdata[52]
port 246 nsew signal input
rlabel metal3 s 0 144304 800 144424 6 dma_hwdata[53]
port 247 nsew signal input
rlabel metal3 s 0 144712 800 144832 6 dma_hwdata[54]
port 248 nsew signal input
rlabel metal3 s 0 145120 800 145240 6 dma_hwdata[55]
port 249 nsew signal input
rlabel metal3 s 0 145392 800 145512 6 dma_hwdata[56]
port 250 nsew signal input
rlabel metal3 s 0 145800 800 145920 6 dma_hwdata[57]
port 251 nsew signal input
rlabel metal3 s 0 146208 800 146328 6 dma_hwdata[58]
port 252 nsew signal input
rlabel metal3 s 0 146480 800 146600 6 dma_hwdata[59]
port 253 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 dma_hwdata[5]
port 254 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 dma_hwdata[60]
port 255 nsew signal input
rlabel metal3 s 0 147160 800 147280 6 dma_hwdata[61]
port 256 nsew signal input
rlabel metal3 s 0 147568 800 147688 6 dma_hwdata[62]
port 257 nsew signal input
rlabel metal3 s 0 147976 800 148096 6 dma_hwdata[63]
port 258 nsew signal input
rlabel metal3 s 0 127576 800 127696 6 dma_hwdata[6]
port 259 nsew signal input
rlabel metal3 s 0 127984 800 128104 6 dma_hwdata[7]
port 260 nsew signal input
rlabel metal3 s 0 128256 800 128376 6 dma_hwdata[8]
port 261 nsew signal input
rlabel metal3 s 0 128664 800 128784 6 dma_hwdata[9]
port 262 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 dma_hwrite
port 263 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 extintsrc_req[0]
port 264 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 extintsrc_req[10]
port 265 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 extintsrc_req[11]
port 266 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 extintsrc_req[12]
port 267 nsew signal input
rlabel metal3 s 0 39312 800 39432 6 extintsrc_req[13]
port 268 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 extintsrc_req[14]
port 269 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 extintsrc_req[15]
port 270 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 extintsrc_req[16]
port 271 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 extintsrc_req[17]
port 272 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 extintsrc_req[18]
port 273 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 extintsrc_req[19]
port 274 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 extintsrc_req[1]
port 275 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 extintsrc_req[20]
port 276 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 extintsrc_req[21]
port 277 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 extintsrc_req[22]
port 278 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 extintsrc_req[23]
port 279 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 extintsrc_req[24]
port 280 nsew signal input
rlabel metal3 s 0 43664 800 43784 6 extintsrc_req[25]
port 281 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 extintsrc_req[26]
port 282 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 extintsrc_req[27]
port 283 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 extintsrc_req[28]
port 284 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 extintsrc_req[29]
port 285 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 extintsrc_req[2]
port 286 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 extintsrc_req[30]
port 287 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 extintsrc_req[3]
port 288 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 extintsrc_req[4]
port 289 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 extintsrc_req[5]
port 290 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 extintsrc_req[6]
port 291 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 extintsrc_req[7]
port 292 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 extintsrc_req[8]
port 293 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 extintsrc_req[9]
port 294 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 haddr[0]
port 295 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 haddr[10]
port 296 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 haddr[11]
port 297 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 haddr[12]
port 298 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 haddr[13]
port 299 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 haddr[14]
port 300 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 haddr[15]
port 301 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 haddr[16]
port 302 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 haddr[17]
port 303 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 haddr[18]
port 304 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 haddr[19]
port 305 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 haddr[1]
port 306 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 haddr[20]
port 307 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 haddr[21]
port 308 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 haddr[22]
port 309 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 haddr[23]
port 310 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 haddr[24]
port 311 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 haddr[25]
port 312 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 haddr[26]
port 313 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 haddr[27]
port 314 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 haddr[28]
port 315 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 haddr[29]
port 316 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 haddr[2]
port 317 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 haddr[30]
port 318 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 haddr[31]
port 319 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 haddr[3]
port 320 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 haddr[4]
port 321 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 haddr[5]
port 322 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 haddr[6]
port 323 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 haddr[7]
port 324 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 haddr[8]
port 325 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 haddr[9]
port 326 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 hburst[0]
port 327 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 hburst[1]
port 328 nsew signal output
rlabel metal3 s 0 28976 800 29096 6 hburst[2]
port 329 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 hmastlock
port 330 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 hprot[0]
port 331 nsew signal output
rlabel metal3 s 0 30064 800 30184 6 hprot[1]
port 332 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 hprot[2]
port 333 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 hprot[3]
port 334 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 hrdata[0]
port 335 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 hrdata[10]
port 336 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 hrdata[11]
port 337 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 hrdata[12]
port 338 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 hrdata[13]
port 339 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 hrdata[14]
port 340 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 hrdata[15]
port 341 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 hrdata[16]
port 342 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 hrdata[17]
port 343 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 hrdata[18]
port 344 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 hrdata[19]
port 345 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 hrdata[1]
port 346 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 hrdata[20]
port 347 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 hrdata[21]
port 348 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 hrdata[22]
port 349 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 hrdata[23]
port 350 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 hrdata[24]
port 351 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 hrdata[25]
port 352 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 hrdata[26]
port 353 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 hrdata[27]
port 354 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 hrdata[28]
port 355 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 hrdata[29]
port 356 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 hrdata[2]
port 357 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 hrdata[30]
port 358 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 hrdata[31]
port 359 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 hrdata[32]
port 360 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 hrdata[33]
port 361 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 hrdata[34]
port 362 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 hrdata[35]
port 363 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 hrdata[36]
port 364 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 hrdata[37]
port 365 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 hrdata[38]
port 366 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 hrdata[39]
port 367 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 hrdata[3]
port 368 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 hrdata[40]
port 369 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 hrdata[41]
port 370 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 hrdata[42]
port 371 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 hrdata[43]
port 372 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 hrdata[44]
port 373 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 hrdata[45]
port 374 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 hrdata[46]
port 375 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 hrdata[47]
port 376 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 hrdata[48]
port 377 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 hrdata[49]
port 378 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 hrdata[4]
port 379 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 hrdata[50]
port 380 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 hrdata[51]
port 381 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 hrdata[52]
port 382 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 hrdata[53]
port 383 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 hrdata[54]
port 384 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 hrdata[55]
port 385 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 hrdata[56]
port 386 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 hrdata[57]
port 387 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 hrdata[58]
port 388 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 hrdata[59]
port 389 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 hrdata[5]
port 390 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 hrdata[60]
port 391 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 hrdata[61]
port 392 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 hrdata[62]
port 393 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 hrdata[63]
port 394 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 hrdata[6]
port 395 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 hrdata[7]
port 396 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 hrdata[8]
port 397 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 hrdata[9]
port 398 nsew signal input
rlabel metal3 s 0 824 800 944 6 hready
port 399 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 hresp
port 400 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 hsize[0]
port 401 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 hsize[1]
port 402 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 hsize[2]
port 403 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 htrans[0]
port 404 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 htrans[1]
port 405 nsew signal output
rlabel metal3 s 0 144 800 264 6 hwrite
port 406 nsew signal output
rlabel metal3 s 0 260040 800 260160 6 i_cpu_halt_req
port 407 nsew signal input
rlabel metal3 s 0 261536 800 261656 6 i_cpu_run_req
port 408 nsew signal input
rlabel metal3 s 0 207952 800 208072 6 ic_data_ext_in_pkt[0]
port 409 nsew signal input
rlabel metal3 s 0 211488 800 211608 6 ic_data_ext_in_pkt[10]
port 410 nsew signal input
rlabel metal3 s 0 211896 800 212016 6 ic_data_ext_in_pkt[11]
port 411 nsew signal input
rlabel metal3 s 0 212168 800 212288 6 ic_data_ext_in_pkt[12]
port 412 nsew signal input
rlabel metal3 s 0 212576 800 212696 6 ic_data_ext_in_pkt[13]
port 413 nsew signal input
rlabel metal3 s 0 212984 800 213104 6 ic_data_ext_in_pkt[14]
port 414 nsew signal input
rlabel metal3 s 0 213256 800 213376 6 ic_data_ext_in_pkt[15]
port 415 nsew signal input
rlabel metal3 s 0 213664 800 213784 6 ic_data_ext_in_pkt[16]
port 416 nsew signal input
rlabel metal3 s 0 214072 800 214192 6 ic_data_ext_in_pkt[17]
port 417 nsew signal input
rlabel metal3 s 0 214344 800 214464 6 ic_data_ext_in_pkt[18]
port 418 nsew signal input
rlabel metal3 s 0 214752 800 214872 6 ic_data_ext_in_pkt[19]
port 419 nsew signal input
rlabel metal3 s 0 208360 800 208480 6 ic_data_ext_in_pkt[1]
port 420 nsew signal input
rlabel metal3 s 0 215024 800 215144 6 ic_data_ext_in_pkt[20]
port 421 nsew signal input
rlabel metal3 s 0 215432 800 215552 6 ic_data_ext_in_pkt[21]
port 422 nsew signal input
rlabel metal3 s 0 215840 800 215960 6 ic_data_ext_in_pkt[22]
port 423 nsew signal input
rlabel metal3 s 0 216112 800 216232 6 ic_data_ext_in_pkt[23]
port 424 nsew signal input
rlabel metal3 s 0 216520 800 216640 6 ic_data_ext_in_pkt[24]
port 425 nsew signal input
rlabel metal3 s 0 216928 800 217048 6 ic_data_ext_in_pkt[25]
port 426 nsew signal input
rlabel metal3 s 0 217200 800 217320 6 ic_data_ext_in_pkt[26]
port 427 nsew signal input
rlabel metal3 s 0 217608 800 217728 6 ic_data_ext_in_pkt[27]
port 428 nsew signal input
rlabel metal3 s 0 217880 800 218000 6 ic_data_ext_in_pkt[28]
port 429 nsew signal input
rlabel metal3 s 0 218288 800 218408 6 ic_data_ext_in_pkt[29]
port 430 nsew signal input
rlabel metal3 s 0 208632 800 208752 6 ic_data_ext_in_pkt[2]
port 431 nsew signal input
rlabel metal3 s 0 218696 800 218816 6 ic_data_ext_in_pkt[30]
port 432 nsew signal input
rlabel metal3 s 0 218968 800 219088 6 ic_data_ext_in_pkt[31]
port 433 nsew signal input
rlabel metal3 s 0 219376 800 219496 6 ic_data_ext_in_pkt[32]
port 434 nsew signal input
rlabel metal3 s 0 219784 800 219904 6 ic_data_ext_in_pkt[33]
port 435 nsew signal input
rlabel metal3 s 0 220056 800 220176 6 ic_data_ext_in_pkt[34]
port 436 nsew signal input
rlabel metal3 s 0 220464 800 220584 6 ic_data_ext_in_pkt[35]
port 437 nsew signal input
rlabel metal3 s 0 220736 800 220856 6 ic_data_ext_in_pkt[36]
port 438 nsew signal input
rlabel metal3 s 0 221144 800 221264 6 ic_data_ext_in_pkt[37]
port 439 nsew signal input
rlabel metal3 s 0 221552 800 221672 6 ic_data_ext_in_pkt[38]
port 440 nsew signal input
rlabel metal3 s 0 221824 800 221944 6 ic_data_ext_in_pkt[39]
port 441 nsew signal input
rlabel metal3 s 0 209040 800 209160 6 ic_data_ext_in_pkt[3]
port 442 nsew signal input
rlabel metal3 s 0 222232 800 222352 6 ic_data_ext_in_pkt[40]
port 443 nsew signal input
rlabel metal3 s 0 222640 800 222760 6 ic_data_ext_in_pkt[41]
port 444 nsew signal input
rlabel metal3 s 0 222912 800 223032 6 ic_data_ext_in_pkt[42]
port 445 nsew signal input
rlabel metal3 s 0 223320 800 223440 6 ic_data_ext_in_pkt[43]
port 446 nsew signal input
rlabel metal3 s 0 223592 800 223712 6 ic_data_ext_in_pkt[44]
port 447 nsew signal input
rlabel metal3 s 0 224000 800 224120 6 ic_data_ext_in_pkt[45]
port 448 nsew signal input
rlabel metal3 s 0 224408 800 224528 6 ic_data_ext_in_pkt[46]
port 449 nsew signal input
rlabel metal3 s 0 224680 800 224800 6 ic_data_ext_in_pkt[47]
port 450 nsew signal input
rlabel metal3 s 0 209312 800 209432 6 ic_data_ext_in_pkt[4]
port 451 nsew signal input
rlabel metal3 s 0 209720 800 209840 6 ic_data_ext_in_pkt[5]
port 452 nsew signal input
rlabel metal3 s 0 210128 800 210248 6 ic_data_ext_in_pkt[6]
port 453 nsew signal input
rlabel metal3 s 0 210400 800 210520 6 ic_data_ext_in_pkt[7]
port 454 nsew signal input
rlabel metal3 s 0 210808 800 210928 6 ic_data_ext_in_pkt[8]
port 455 nsew signal input
rlabel metal3 s 0 211216 800 211336 6 ic_data_ext_in_pkt[9]
port 456 nsew signal input
rlabel metal3 s 0 225088 800 225208 6 ic_tag_ext_in_pkt[0]
port 457 nsew signal input
rlabel metal3 s 0 228624 800 228744 6 ic_tag_ext_in_pkt[10]
port 458 nsew signal input
rlabel metal3 s 0 229032 800 229152 6 ic_tag_ext_in_pkt[11]
port 459 nsew signal input
rlabel metal3 s 0 229440 800 229560 6 ic_tag_ext_in_pkt[12]
port 460 nsew signal input
rlabel metal3 s 0 229712 800 229832 6 ic_tag_ext_in_pkt[13]
port 461 nsew signal input
rlabel metal3 s 0 230120 800 230240 6 ic_tag_ext_in_pkt[14]
port 462 nsew signal input
rlabel metal3 s 0 230392 800 230512 6 ic_tag_ext_in_pkt[15]
port 463 nsew signal input
rlabel metal3 s 0 230800 800 230920 6 ic_tag_ext_in_pkt[16]
port 464 nsew signal input
rlabel metal3 s 0 231208 800 231328 6 ic_tag_ext_in_pkt[17]
port 465 nsew signal input
rlabel metal3 s 0 231480 800 231600 6 ic_tag_ext_in_pkt[18]
port 466 nsew signal input
rlabel metal3 s 0 231888 800 232008 6 ic_tag_ext_in_pkt[19]
port 467 nsew signal input
rlabel metal3 s 0 225496 800 225616 6 ic_tag_ext_in_pkt[1]
port 468 nsew signal input
rlabel metal3 s 0 232296 800 232416 6 ic_tag_ext_in_pkt[20]
port 469 nsew signal input
rlabel metal3 s 0 232568 800 232688 6 ic_tag_ext_in_pkt[21]
port 470 nsew signal input
rlabel metal3 s 0 232976 800 233096 6 ic_tag_ext_in_pkt[22]
port 471 nsew signal input
rlabel metal3 s 0 233248 800 233368 6 ic_tag_ext_in_pkt[23]
port 472 nsew signal input
rlabel metal3 s 0 225768 800 225888 6 ic_tag_ext_in_pkt[2]
port 473 nsew signal input
rlabel metal3 s 0 226176 800 226296 6 ic_tag_ext_in_pkt[3]
port 474 nsew signal input
rlabel metal3 s 0 226584 800 226704 6 ic_tag_ext_in_pkt[4]
port 475 nsew signal input
rlabel metal3 s 0 226856 800 226976 6 ic_tag_ext_in_pkt[5]
port 476 nsew signal input
rlabel metal3 s 0 227264 800 227384 6 ic_tag_ext_in_pkt[6]
port 477 nsew signal input
rlabel metal3 s 0 227536 800 227656 6 ic_tag_ext_in_pkt[7]
port 478 nsew signal input
rlabel metal3 s 0 227944 800 228064 6 ic_tag_ext_in_pkt[8]
port 479 nsew signal input
rlabel metal3 s 0 228352 800 228472 6 ic_tag_ext_in_pkt[9]
port 480 nsew signal input
rlabel metal3 s 0 190816 800 190936 6 iccm_ext_in_pkt[0]
port 481 nsew signal input
rlabel metal3 s 0 194352 800 194472 6 iccm_ext_in_pkt[10]
port 482 nsew signal input
rlabel metal3 s 0 194760 800 194880 6 iccm_ext_in_pkt[11]
port 483 nsew signal input
rlabel metal3 s 0 195032 800 195152 6 iccm_ext_in_pkt[12]
port 484 nsew signal input
rlabel metal3 s 0 195440 800 195560 6 iccm_ext_in_pkt[13]
port 485 nsew signal input
rlabel metal3 s 0 195848 800 195968 6 iccm_ext_in_pkt[14]
port 486 nsew signal input
rlabel metal3 s 0 196120 800 196240 6 iccm_ext_in_pkt[15]
port 487 nsew signal input
rlabel metal3 s 0 196528 800 196648 6 iccm_ext_in_pkt[16]
port 488 nsew signal input
rlabel metal3 s 0 196936 800 197056 6 iccm_ext_in_pkt[17]
port 489 nsew signal input
rlabel metal3 s 0 197208 800 197328 6 iccm_ext_in_pkt[18]
port 490 nsew signal input
rlabel metal3 s 0 197616 800 197736 6 iccm_ext_in_pkt[19]
port 491 nsew signal input
rlabel metal3 s 0 191224 800 191344 6 iccm_ext_in_pkt[1]
port 492 nsew signal input
rlabel metal3 s 0 197888 800 198008 6 iccm_ext_in_pkt[20]
port 493 nsew signal input
rlabel metal3 s 0 198296 800 198416 6 iccm_ext_in_pkt[21]
port 494 nsew signal input
rlabel metal3 s 0 198704 800 198824 6 iccm_ext_in_pkt[22]
port 495 nsew signal input
rlabel metal3 s 0 198976 800 199096 6 iccm_ext_in_pkt[23]
port 496 nsew signal input
rlabel metal3 s 0 199384 800 199504 6 iccm_ext_in_pkt[24]
port 497 nsew signal input
rlabel metal3 s 0 199792 800 199912 6 iccm_ext_in_pkt[25]
port 498 nsew signal input
rlabel metal3 s 0 200064 800 200184 6 iccm_ext_in_pkt[26]
port 499 nsew signal input
rlabel metal3 s 0 200472 800 200592 6 iccm_ext_in_pkt[27]
port 500 nsew signal input
rlabel metal3 s 0 200744 800 200864 6 iccm_ext_in_pkt[28]
port 501 nsew signal input
rlabel metal3 s 0 201152 800 201272 6 iccm_ext_in_pkt[29]
port 502 nsew signal input
rlabel metal3 s 0 191496 800 191616 6 iccm_ext_in_pkt[2]
port 503 nsew signal input
rlabel metal3 s 0 201560 800 201680 6 iccm_ext_in_pkt[30]
port 504 nsew signal input
rlabel metal3 s 0 201832 800 201952 6 iccm_ext_in_pkt[31]
port 505 nsew signal input
rlabel metal3 s 0 202240 800 202360 6 iccm_ext_in_pkt[32]
port 506 nsew signal input
rlabel metal3 s 0 202648 800 202768 6 iccm_ext_in_pkt[33]
port 507 nsew signal input
rlabel metal3 s 0 202920 800 203040 6 iccm_ext_in_pkt[34]
port 508 nsew signal input
rlabel metal3 s 0 203328 800 203448 6 iccm_ext_in_pkt[35]
port 509 nsew signal input
rlabel metal3 s 0 203600 800 203720 6 iccm_ext_in_pkt[36]
port 510 nsew signal input
rlabel metal3 s 0 204008 800 204128 6 iccm_ext_in_pkt[37]
port 511 nsew signal input
rlabel metal3 s 0 204416 800 204536 6 iccm_ext_in_pkt[38]
port 512 nsew signal input
rlabel metal3 s 0 204688 800 204808 6 iccm_ext_in_pkt[39]
port 513 nsew signal input
rlabel metal3 s 0 191904 800 192024 6 iccm_ext_in_pkt[3]
port 514 nsew signal input
rlabel metal3 s 0 205096 800 205216 6 iccm_ext_in_pkt[40]
port 515 nsew signal input
rlabel metal3 s 0 205504 800 205624 6 iccm_ext_in_pkt[41]
port 516 nsew signal input
rlabel metal3 s 0 205776 800 205896 6 iccm_ext_in_pkt[42]
port 517 nsew signal input
rlabel metal3 s 0 206184 800 206304 6 iccm_ext_in_pkt[43]
port 518 nsew signal input
rlabel metal3 s 0 206456 800 206576 6 iccm_ext_in_pkt[44]
port 519 nsew signal input
rlabel metal3 s 0 206864 800 206984 6 iccm_ext_in_pkt[45]
port 520 nsew signal input
rlabel metal3 s 0 207272 800 207392 6 iccm_ext_in_pkt[46]
port 521 nsew signal input
rlabel metal3 s 0 207544 800 207664 6 iccm_ext_in_pkt[47]
port 522 nsew signal input
rlabel metal3 s 0 192176 800 192296 6 iccm_ext_in_pkt[4]
port 523 nsew signal input
rlabel metal3 s 0 192584 800 192704 6 iccm_ext_in_pkt[5]
port 524 nsew signal input
rlabel metal3 s 0 192992 800 193112 6 iccm_ext_in_pkt[6]
port 525 nsew signal input
rlabel metal3 s 0 193264 800 193384 6 iccm_ext_in_pkt[7]
port 526 nsew signal input
rlabel metal3 s 0 193672 800 193792 6 iccm_ext_in_pkt[8]
port 527 nsew signal input
rlabel metal3 s 0 194080 800 194200 6 iccm_ext_in_pkt[9]
port 528 nsew signal input
rlabel metal3 s 0 172592 800 172712 6 ifu_bus_clk_en
port 529 nsew signal input
rlabel metal3 s 0 236920 800 237040 6 jtag_id[0]
port 530 nsew signal input
rlabel metal3 s 0 240456 800 240576 6 jtag_id[10]
port 531 nsew signal input
rlabel metal3 s 0 240864 800 240984 6 jtag_id[11]
port 532 nsew signal input
rlabel metal3 s 0 241136 800 241256 6 jtag_id[12]
port 533 nsew signal input
rlabel metal3 s 0 241544 800 241664 6 jtag_id[13]
port 534 nsew signal input
rlabel metal3 s 0 241816 800 241936 6 jtag_id[14]
port 535 nsew signal input
rlabel metal3 s 0 242224 800 242344 6 jtag_id[15]
port 536 nsew signal input
rlabel metal3 s 0 242632 800 242752 6 jtag_id[16]
port 537 nsew signal input
rlabel metal3 s 0 242904 800 243024 6 jtag_id[17]
port 538 nsew signal input
rlabel metal3 s 0 243312 800 243432 6 jtag_id[18]
port 539 nsew signal input
rlabel metal3 s 0 243720 800 243840 6 jtag_id[19]
port 540 nsew signal input
rlabel metal3 s 0 237192 800 237312 6 jtag_id[1]
port 541 nsew signal input
rlabel metal3 s 0 243992 800 244112 6 jtag_id[20]
port 542 nsew signal input
rlabel metal3 s 0 244400 800 244520 6 jtag_id[21]
port 543 nsew signal input
rlabel metal3 s 0 244672 800 244792 6 jtag_id[22]
port 544 nsew signal input
rlabel metal3 s 0 245080 800 245200 6 jtag_id[23]
port 545 nsew signal input
rlabel metal3 s 0 245488 800 245608 6 jtag_id[24]
port 546 nsew signal input
rlabel metal3 s 0 245760 800 245880 6 jtag_id[25]
port 547 nsew signal input
rlabel metal3 s 0 246168 800 246288 6 jtag_id[26]
port 548 nsew signal input
rlabel metal3 s 0 246576 800 246696 6 jtag_id[27]
port 549 nsew signal input
rlabel metal3 s 0 246848 800 246968 6 jtag_id[28]
port 550 nsew signal input
rlabel metal3 s 0 247256 800 247376 6 jtag_id[29]
port 551 nsew signal input
rlabel metal3 s 0 237600 800 237720 6 jtag_id[2]
port 552 nsew signal input
rlabel metal3 s 0 247528 800 247648 6 jtag_id[30]
port 553 nsew signal input
rlabel metal3 s 0 238008 800 238128 6 jtag_id[3]
port 554 nsew signal input
rlabel metal3 s 0 238280 800 238400 6 jtag_id[4]
port 555 nsew signal input
rlabel metal3 s 0 238688 800 238808 6 jtag_id[5]
port 556 nsew signal input
rlabel metal3 s 0 238960 800 239080 6 jtag_id[6]
port 557 nsew signal input
rlabel metal3 s 0 239368 800 239488 6 jtag_id[7]
port 558 nsew signal input
rlabel metal3 s 0 239776 800 239896 6 jtag_id[8]
port 559 nsew signal input
rlabel metal3 s 0 240048 800 240168 6 jtag_id[9]
port 560 nsew signal input
rlabel metal3 s 0 235152 800 235272 6 jtag_tck
port 561 nsew signal input
rlabel metal3 s 0 235832 800 235952 6 jtag_tdi
port 562 nsew signal input
rlabel metal3 s 0 236512 800 236632 6 jtag_tdo
port 563 nsew signal output
rlabel metal3 s 0 235424 800 235544 6 jtag_tms
port 564 nsew signal input
rlabel metal3 s 0 236104 800 236224 6 jtag_trst_n
port 565 nsew signal input
rlabel metal3 s 0 172184 800 172304 6 lsu_bus_clk_en
port 566 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 lsu_haddr[0]
port 567 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 lsu_haddr[10]
port 568 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 lsu_haddr[11]
port 569 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 lsu_haddr[12]
port 570 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 lsu_haddr[13]
port 571 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 lsu_haddr[14]
port 572 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 lsu_haddr[15]
port 573 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 lsu_haddr[16]
port 574 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 lsu_haddr[17]
port 575 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 lsu_haddr[18]
port 576 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 lsu_haddr[19]
port 577 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 lsu_haddr[1]
port 578 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 lsu_haddr[20]
port 579 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 lsu_haddr[21]
port 580 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 lsu_haddr[22]
port 581 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 lsu_haddr[23]
port 582 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 lsu_haddr[24]
port 583 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 lsu_haddr[25]
port 584 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 lsu_haddr[26]
port 585 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 lsu_haddr[27]
port 586 nsew signal output
rlabel metal2 s 68558 0 68614 800 6 lsu_haddr[28]
port 587 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 lsu_haddr[29]
port 588 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 lsu_haddr[2]
port 589 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 lsu_haddr[30]
port 590 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 lsu_haddr[31]
port 591 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 lsu_haddr[3]
port 592 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 lsu_haddr[4]
port 593 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 lsu_haddr[5]
port 594 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 lsu_haddr[6]
port 595 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 lsu_haddr[7]
port 596 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 lsu_haddr[8]
port 597 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 lsu_haddr[9]
port 598 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 lsu_hburst[0]
port 599 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 lsu_hburst[1]
port 600 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 lsu_hburst[2]
port 601 nsew signal output
rlabel metal3 s 0 32240 800 32360 6 lsu_hmastlock
port 602 nsew signal output
rlabel metal3 s 0 32512 800 32632 6 lsu_hprot[0]
port 603 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 lsu_hprot[1]
port 604 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 lsu_hprot[2]
port 605 nsew signal output
rlabel metal3 s 0 33600 800 33720 6 lsu_hprot[3]
port 606 nsew signal output
rlabel metal2 s 142066 0 142122 800 6 lsu_hrdata[0]
port 607 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 lsu_hrdata[10]
port 608 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 lsu_hrdata[11]
port 609 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 lsu_hrdata[12]
port 610 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 lsu_hrdata[13]
port 611 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 lsu_hrdata[14]
port 612 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 lsu_hrdata[15]
port 613 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 lsu_hrdata[16]
port 614 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 lsu_hrdata[17]
port 615 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 lsu_hrdata[18]
port 616 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 lsu_hrdata[19]
port 617 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 lsu_hrdata[1]
port 618 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 lsu_hrdata[20]
port 619 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 lsu_hrdata[21]
port 620 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 lsu_hrdata[22]
port 621 nsew signal input
rlabel metal2 s 166906 0 166962 800 6 lsu_hrdata[23]
port 622 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 lsu_hrdata[24]
port 623 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 lsu_hrdata[25]
port 624 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 lsu_hrdata[26]
port 625 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 lsu_hrdata[27]
port 626 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 lsu_hrdata[28]
port 627 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 lsu_hrdata[29]
port 628 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 lsu_hrdata[2]
port 629 nsew signal input
rlabel metal2 s 174450 0 174506 800 6 lsu_hrdata[30]
port 630 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 lsu_hrdata[31]
port 631 nsew signal input
rlabel metal2 s 176658 0 176714 800 6 lsu_hrdata[32]
port 632 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 lsu_hrdata[33]
port 633 nsew signal input
rlabel metal2 s 178774 0 178830 800 6 lsu_hrdata[34]
port 634 nsew signal input
rlabel metal2 s 179878 0 179934 800 6 lsu_hrdata[35]
port 635 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 lsu_hrdata[36]
port 636 nsew signal input
rlabel metal2 s 181994 0 182050 800 6 lsu_hrdata[37]
port 637 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 lsu_hrdata[38]
port 638 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 lsu_hrdata[39]
port 639 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 lsu_hrdata[3]
port 640 nsew signal input
rlabel metal2 s 185306 0 185362 800 6 lsu_hrdata[40]
port 641 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 lsu_hrdata[41]
port 642 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 lsu_hrdata[42]
port 643 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 lsu_hrdata[43]
port 644 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 lsu_hrdata[44]
port 645 nsew signal input
rlabel metal2 s 190642 0 190698 800 6 lsu_hrdata[45]
port 646 nsew signal input
rlabel metal2 s 191746 0 191802 800 6 lsu_hrdata[46]
port 647 nsew signal input
rlabel metal2 s 192850 0 192906 800 6 lsu_hrdata[47]
port 648 nsew signal input
rlabel metal2 s 193954 0 194010 800 6 lsu_hrdata[48]
port 649 nsew signal input
rlabel metal2 s 194966 0 195022 800 6 lsu_hrdata[49]
port 650 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 lsu_hrdata[4]
port 651 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 lsu_hrdata[50]
port 652 nsew signal input
rlabel metal2 s 197174 0 197230 800 6 lsu_hrdata[51]
port 653 nsew signal input
rlabel metal2 s 198278 0 198334 800 6 lsu_hrdata[52]
port 654 nsew signal input
rlabel metal2 s 199290 0 199346 800 6 lsu_hrdata[53]
port 655 nsew signal input
rlabel metal2 s 200394 0 200450 800 6 lsu_hrdata[54]
port 656 nsew signal input
rlabel metal2 s 201498 0 201554 800 6 lsu_hrdata[55]
port 657 nsew signal input
rlabel metal2 s 202602 0 202658 800 6 lsu_hrdata[56]
port 658 nsew signal input
rlabel metal2 s 203614 0 203670 800 6 lsu_hrdata[57]
port 659 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 lsu_hrdata[58]
port 660 nsew signal input
rlabel metal2 s 205822 0 205878 800 6 lsu_hrdata[59]
port 661 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 lsu_hrdata[5]
port 662 nsew signal input
rlabel metal2 s 206926 0 206982 800 6 lsu_hrdata[60]
port 663 nsew signal input
rlabel metal2 s 207938 0 207994 800 6 lsu_hrdata[61]
port 664 nsew signal input
rlabel metal2 s 209042 0 209098 800 6 lsu_hrdata[62]
port 665 nsew signal input
rlabel metal2 s 210146 0 210202 800 6 lsu_hrdata[63]
port 666 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 lsu_hrdata[6]
port 667 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 lsu_hrdata[7]
port 668 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 lsu_hrdata[8]
port 669 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 lsu_hrdata[9]
port 670 nsew signal input
rlabel metal3 s 0 1096 800 1216 6 lsu_hready
port 671 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 lsu_hresp
port 672 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 lsu_hsize[0]
port 673 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 lsu_hsize[1]
port 674 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 lsu_hsize[2]
port 675 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 lsu_htrans[0]
port 676 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 lsu_htrans[1]
port 677 nsew signal output
rlabel metal2 s 211250 0 211306 800 6 lsu_hwdata[0]
port 678 nsew signal output
rlabel metal2 s 222014 0 222070 800 6 lsu_hwdata[10]
port 679 nsew signal output
rlabel metal2 s 223118 0 223174 800 6 lsu_hwdata[11]
port 680 nsew signal output
rlabel metal2 s 224222 0 224278 800 6 lsu_hwdata[12]
port 681 nsew signal output
rlabel metal2 s 225234 0 225290 800 6 lsu_hwdata[13]
port 682 nsew signal output
rlabel metal2 s 226338 0 226394 800 6 lsu_hwdata[14]
port 683 nsew signal output
rlabel metal2 s 227442 0 227498 800 6 lsu_hwdata[15]
port 684 nsew signal output
rlabel metal2 s 228546 0 228602 800 6 lsu_hwdata[16]
port 685 nsew signal output
rlabel metal2 s 229558 0 229614 800 6 lsu_hwdata[17]
port 686 nsew signal output
rlabel metal2 s 230662 0 230718 800 6 lsu_hwdata[18]
port 687 nsew signal output
rlabel metal2 s 231766 0 231822 800 6 lsu_hwdata[19]
port 688 nsew signal output
rlabel metal2 s 212262 0 212318 800 6 lsu_hwdata[1]
port 689 nsew signal output
rlabel metal2 s 232870 0 232926 800 6 lsu_hwdata[20]
port 690 nsew signal output
rlabel metal2 s 233882 0 233938 800 6 lsu_hwdata[21]
port 691 nsew signal output
rlabel metal2 s 234986 0 235042 800 6 lsu_hwdata[22]
port 692 nsew signal output
rlabel metal2 s 236090 0 236146 800 6 lsu_hwdata[23]
port 693 nsew signal output
rlabel metal2 s 237194 0 237250 800 6 lsu_hwdata[24]
port 694 nsew signal output
rlabel metal2 s 238206 0 238262 800 6 lsu_hwdata[25]
port 695 nsew signal output
rlabel metal2 s 239310 0 239366 800 6 lsu_hwdata[26]
port 696 nsew signal output
rlabel metal2 s 240414 0 240470 800 6 lsu_hwdata[27]
port 697 nsew signal output
rlabel metal2 s 241518 0 241574 800 6 lsu_hwdata[28]
port 698 nsew signal output
rlabel metal2 s 242530 0 242586 800 6 lsu_hwdata[29]
port 699 nsew signal output
rlabel metal2 s 213366 0 213422 800 6 lsu_hwdata[2]
port 700 nsew signal output
rlabel metal2 s 243634 0 243690 800 6 lsu_hwdata[30]
port 701 nsew signal output
rlabel metal2 s 244738 0 244794 800 6 lsu_hwdata[31]
port 702 nsew signal output
rlabel metal2 s 245842 0 245898 800 6 lsu_hwdata[32]
port 703 nsew signal output
rlabel metal2 s 246854 0 246910 800 6 lsu_hwdata[33]
port 704 nsew signal output
rlabel metal2 s 247958 0 248014 800 6 lsu_hwdata[34]
port 705 nsew signal output
rlabel metal2 s 249062 0 249118 800 6 lsu_hwdata[35]
port 706 nsew signal output
rlabel metal2 s 250166 0 250222 800 6 lsu_hwdata[36]
port 707 nsew signal output
rlabel metal2 s 251178 0 251234 800 6 lsu_hwdata[37]
port 708 nsew signal output
rlabel metal2 s 252282 0 252338 800 6 lsu_hwdata[38]
port 709 nsew signal output
rlabel metal2 s 253386 0 253442 800 6 lsu_hwdata[39]
port 710 nsew signal output
rlabel metal2 s 214470 0 214526 800 6 lsu_hwdata[3]
port 711 nsew signal output
rlabel metal2 s 254490 0 254546 800 6 lsu_hwdata[40]
port 712 nsew signal output
rlabel metal2 s 255502 0 255558 800 6 lsu_hwdata[41]
port 713 nsew signal output
rlabel metal2 s 256606 0 256662 800 6 lsu_hwdata[42]
port 714 nsew signal output
rlabel metal2 s 257710 0 257766 800 6 lsu_hwdata[43]
port 715 nsew signal output
rlabel metal2 s 258814 0 258870 800 6 lsu_hwdata[44]
port 716 nsew signal output
rlabel metal2 s 259826 0 259882 800 6 lsu_hwdata[45]
port 717 nsew signal output
rlabel metal2 s 260930 0 260986 800 6 lsu_hwdata[46]
port 718 nsew signal output
rlabel metal2 s 262034 0 262090 800 6 lsu_hwdata[47]
port 719 nsew signal output
rlabel metal2 s 263138 0 263194 800 6 lsu_hwdata[48]
port 720 nsew signal output
rlabel metal2 s 264150 0 264206 800 6 lsu_hwdata[49]
port 721 nsew signal output
rlabel metal2 s 215574 0 215630 800 6 lsu_hwdata[4]
port 722 nsew signal output
rlabel metal2 s 265254 0 265310 800 6 lsu_hwdata[50]
port 723 nsew signal output
rlabel metal2 s 266358 0 266414 800 6 lsu_hwdata[51]
port 724 nsew signal output
rlabel metal2 s 267462 0 267518 800 6 lsu_hwdata[52]
port 725 nsew signal output
rlabel metal2 s 268474 0 268530 800 6 lsu_hwdata[53]
port 726 nsew signal output
rlabel metal2 s 269578 0 269634 800 6 lsu_hwdata[54]
port 727 nsew signal output
rlabel metal2 s 270682 0 270738 800 6 lsu_hwdata[55]
port 728 nsew signal output
rlabel metal2 s 271786 0 271842 800 6 lsu_hwdata[56]
port 729 nsew signal output
rlabel metal2 s 272798 0 272854 800 6 lsu_hwdata[57]
port 730 nsew signal output
rlabel metal2 s 273902 0 273958 800 6 lsu_hwdata[58]
port 731 nsew signal output
rlabel metal2 s 275006 0 275062 800 6 lsu_hwdata[59]
port 732 nsew signal output
rlabel metal2 s 216586 0 216642 800 6 lsu_hwdata[5]
port 733 nsew signal output
rlabel metal2 s 276110 0 276166 800 6 lsu_hwdata[60]
port 734 nsew signal output
rlabel metal2 s 277122 0 277178 800 6 lsu_hwdata[61]
port 735 nsew signal output
rlabel metal2 s 278226 0 278282 800 6 lsu_hwdata[62]
port 736 nsew signal output
rlabel metal2 s 279330 0 279386 800 6 lsu_hwdata[63]
port 737 nsew signal output
rlabel metal2 s 217690 0 217746 800 6 lsu_hwdata[6]
port 738 nsew signal output
rlabel metal2 s 218794 0 218850 800 6 lsu_hwdata[7]
port 739 nsew signal output
rlabel metal2 s 219898 0 219954 800 6 lsu_hwdata[8]
port 740 nsew signal output
rlabel metal2 s 220910 0 220966 800 6 lsu_hwdata[9]
port 741 nsew signal output
rlabel metal3 s 0 416 800 536 6 lsu_hwrite
port 742 nsew signal output
rlabel metal3 s 0 262624 800 262744 6 mbist_mode
port 743 nsew signal input
rlabel metal3 s 0 258952 800 259072 6 mpc_debug_halt_ack
port 744 nsew signal output
rlabel metal3 s 0 258000 800 258120 6 mpc_debug_halt_req
port 745 nsew signal input
rlabel metal3 s 0 259360 800 259480 6 mpc_debug_run_ack
port 746 nsew signal output
rlabel metal3 s 0 258272 800 258392 6 mpc_debug_run_req
port 747 nsew signal input
rlabel metal3 s 0 258680 800 258800 6 mpc_reset_run_req
port 748 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 nmi_int
port 749 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 nmi_vec[0]
port 750 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 nmi_vec[10]
port 751 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 nmi_vec[11]
port 752 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 nmi_vec[12]
port 753 nsew signal input
rlabel metal3 s 0 17552 800 17672 6 nmi_vec[13]
port 754 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 nmi_vec[14]
port 755 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 nmi_vec[15]
port 756 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 nmi_vec[16]
port 757 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 nmi_vec[17]
port 758 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 nmi_vec[18]
port 759 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 nmi_vec[19]
port 760 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 nmi_vec[1]
port 761 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 nmi_vec[20]
port 762 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 nmi_vec[21]
port 763 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 nmi_vec[22]
port 764 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 nmi_vec[23]
port 765 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 nmi_vec[24]
port 766 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 nmi_vec[25]
port 767 nsew signal input
rlabel metal3 s 0 22176 800 22296 6 nmi_vec[26]
port 768 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 nmi_vec[27]
port 769 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 nmi_vec[28]
port 770 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 nmi_vec[29]
port 771 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 nmi_vec[2]
port 772 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 nmi_vec[30]
port 773 nsew signal input
rlabel metal3 s 0 14016 800 14136 6 nmi_vec[3]
port 774 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 nmi_vec[4]
port 775 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 nmi_vec[5]
port 776 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 nmi_vec[6]
port 777 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 nmi_vec[7]
port 778 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 nmi_vec[8]
port 779 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 nmi_vec[9]
port 780 nsew signal input
rlabel metal3 s 0 260448 800 260568 6 o_cpu_halt_ack
port 781 nsew signal output
rlabel metal3 s 0 260856 800 260976 6 o_cpu_halt_status
port 782 nsew signal output
rlabel metal3 s 0 261808 800 261928 6 o_cpu_run_ack
port 783 nsew signal output
rlabel metal3 s 0 261128 800 261248 6 o_debug_mode_status
port 784 nsew signal output
rlabel metal2 s 1490 0 1546 800 6 rst_l
port 785 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 rst_vec[0]
port 786 nsew signal input
rlabel metal3 s 0 5040 800 5160 6 rst_vec[10]
port 787 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 rst_vec[11]
port 788 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 rst_vec[12]
port 789 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 rst_vec[13]
port 790 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 rst_vec[14]
port 791 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 rst_vec[15]
port 792 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 rst_vec[16]
port 793 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 rst_vec[17]
port 794 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 rst_vec[18]
port 795 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 rst_vec[19]
port 796 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 rst_vec[1]
port 797 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 rst_vec[20]
port 798 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 rst_vec[21]
port 799 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 rst_vec[22]
port 800 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 rst_vec[23]
port 801 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 rst_vec[24]
port 802 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 rst_vec[25]
port 803 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 rst_vec[26]
port 804 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 rst_vec[27]
port 805 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 rst_vec[28]
port 806 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 rst_vec[29]
port 807 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 rst_vec[2]
port 808 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 rst_vec[30]
port 809 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 rst_vec[3]
port 810 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 rst_vec[4]
port 811 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 rst_vec[5]
port 812 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 rst_vec[6]
port 813 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 rst_vec[7]
port 814 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 rst_vec[8]
port 815 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 rst_vec[9]
port 816 nsew signal input
rlabel metal3 s 0 45840 800 45960 6 sb_haddr[0]
port 817 nsew signal output
rlabel metal3 s 0 49376 800 49496 6 sb_haddr[10]
port 818 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 sb_haddr[11]
port 819 nsew signal output
rlabel metal3 s 0 50056 800 50176 6 sb_haddr[12]
port 820 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 sb_haddr[13]
port 821 nsew signal output
rlabel metal3 s 0 50736 800 50856 6 sb_haddr[14]
port 822 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 sb_haddr[15]
port 823 nsew signal output
rlabel metal3 s 0 51552 800 51672 6 sb_haddr[16]
port 824 nsew signal output
rlabel metal3 s 0 51824 800 51944 6 sb_haddr[17]
port 825 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 sb_haddr[18]
port 826 nsew signal output
rlabel metal3 s 0 52640 800 52760 6 sb_haddr[19]
port 827 nsew signal output
rlabel metal3 s 0 46112 800 46232 6 sb_haddr[1]
port 828 nsew signal output
rlabel metal3 s 0 52912 800 53032 6 sb_haddr[20]
port 829 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 sb_haddr[21]
port 830 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 sb_haddr[22]
port 831 nsew signal output
rlabel metal3 s 0 54000 800 54120 6 sb_haddr[23]
port 832 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 sb_haddr[24]
port 833 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 sb_haddr[25]
port 834 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 sb_haddr[26]
port 835 nsew signal output
rlabel metal3 s 0 55496 800 55616 6 sb_haddr[27]
port 836 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 sb_haddr[28]
port 837 nsew signal output
rlabel metal3 s 0 56176 800 56296 6 sb_haddr[29]
port 838 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 sb_haddr[2]
port 839 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 sb_haddr[30]
port 840 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 sb_haddr[31]
port 841 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 sb_haddr[3]
port 842 nsew signal output
rlabel metal3 s 0 47200 800 47320 6 sb_haddr[4]
port 843 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 sb_haddr[5]
port 844 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 sb_haddr[6]
port 845 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 sb_haddr[7]
port 846 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 sb_haddr[8]
port 847 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 sb_haddr[9]
port 848 nsew signal output
rlabel metal3 s 0 57264 800 57384 6 sb_hburst[0]
port 849 nsew signal output
rlabel metal3 s 0 57536 800 57656 6 sb_hburst[1]
port 850 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 sb_hburst[2]
port 851 nsew signal output
rlabel metal3 s 0 58352 800 58472 6 sb_hmastlock
port 852 nsew signal output
rlabel metal3 s 0 58624 800 58744 6 sb_hprot[0]
port 853 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 sb_hprot[1]
port 854 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 sb_hprot[2]
port 855 nsew signal output
rlabel metal3 s 0 59712 800 59832 6 sb_hprot[3]
port 856 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 sb_hrdata[0]
port 857 nsew signal input
rlabel metal3 s 0 88680 800 88800 6 sb_hrdata[10]
port 858 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 sb_hrdata[11]
port 859 nsew signal input
rlabel metal3 s 0 89360 800 89480 6 sb_hrdata[12]
port 860 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 sb_hrdata[13]
port 861 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 sb_hrdata[14]
port 862 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 sb_hrdata[15]
port 863 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 sb_hrdata[16]
port 864 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 sb_hrdata[17]
port 865 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 sb_hrdata[18]
port 866 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 sb_hrdata[19]
port 867 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 sb_hrdata[1]
port 868 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 sb_hrdata[20]
port 869 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 sb_hrdata[21]
port 870 nsew signal input
rlabel metal3 s 0 92896 800 93016 6 sb_hrdata[22]
port 871 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 sb_hrdata[23]
port 872 nsew signal input
rlabel metal3 s 0 93712 800 93832 6 sb_hrdata[24]
port 873 nsew signal input
rlabel metal3 s 0 93984 800 94104 6 sb_hrdata[25]
port 874 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 sb_hrdata[26]
port 875 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 sb_hrdata[27]
port 876 nsew signal input
rlabel metal3 s 0 95072 800 95192 6 sb_hrdata[28]
port 877 nsew signal input
rlabel metal3 s 0 95480 800 95600 6 sb_hrdata[29]
port 878 nsew signal input
rlabel metal3 s 0 85824 800 85944 6 sb_hrdata[2]
port 879 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 sb_hrdata[30]
port 880 nsew signal input
rlabel metal3 s 0 96160 800 96280 6 sb_hrdata[31]
port 881 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 sb_hrdata[32]
port 882 nsew signal input
rlabel metal3 s 0 96840 800 96960 6 sb_hrdata[33]
port 883 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 sb_hrdata[34]
port 884 nsew signal input
rlabel metal3 s 0 97520 800 97640 6 sb_hrdata[35]
port 885 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 sb_hrdata[36]
port 886 nsew signal input
rlabel metal3 s 0 98336 800 98456 6 sb_hrdata[37]
port 887 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 sb_hrdata[38]
port 888 nsew signal input
rlabel metal3 s 0 99016 800 99136 6 sb_hrdata[39]
port 889 nsew signal input
rlabel metal3 s 0 86096 800 86216 6 sb_hrdata[3]
port 890 nsew signal input
rlabel metal3 s 0 99424 800 99544 6 sb_hrdata[40]
port 891 nsew signal input
rlabel metal3 s 0 99696 800 99816 6 sb_hrdata[41]
port 892 nsew signal input
rlabel metal3 s 0 100104 800 100224 6 sb_hrdata[42]
port 893 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 sb_hrdata[43]
port 894 nsew signal input
rlabel metal3 s 0 100784 800 100904 6 sb_hrdata[44]
port 895 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 sb_hrdata[45]
port 896 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 sb_hrdata[46]
port 897 nsew signal input
rlabel metal3 s 0 101872 800 101992 6 sb_hrdata[47]
port 898 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 sb_hrdata[48]
port 899 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 sb_hrdata[49]
port 900 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 sb_hrdata[4]
port 901 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 sb_hrdata[50]
port 902 nsew signal input
rlabel metal3 s 0 103232 800 103352 6 sb_hrdata[51]
port 903 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 sb_hrdata[52]
port 904 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 sb_hrdata[53]
port 905 nsew signal input
rlabel metal3 s 0 104320 800 104440 6 sb_hrdata[54]
port 906 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 sb_hrdata[55]
port 907 nsew signal input
rlabel metal3 s 0 105136 800 105256 6 sb_hrdata[56]
port 908 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 sb_hrdata[57]
port 909 nsew signal input
rlabel metal3 s 0 105816 800 105936 6 sb_hrdata[58]
port 910 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 sb_hrdata[59]
port 911 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 sb_hrdata[5]
port 912 nsew signal input
rlabel metal3 s 0 106496 800 106616 6 sb_hrdata[60]
port 913 nsew signal input
rlabel metal3 s 0 106904 800 107024 6 sb_hrdata[61]
port 914 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 sb_hrdata[62]
port 915 nsew signal input
rlabel metal3 s 0 107584 800 107704 6 sb_hrdata[63]
port 916 nsew signal input
rlabel metal3 s 0 87184 800 87304 6 sb_hrdata[6]
port 917 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 sb_hrdata[7]
port 918 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 sb_hrdata[8]
port 919 nsew signal input
rlabel metal3 s 0 88272 800 88392 6 sb_hrdata[9]
port 920 nsew signal input
rlabel metal3 s 0 107992 800 108112 6 sb_hready
port 921 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 sb_hresp
port 922 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 sb_hsize[0]
port 923 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 sb_hsize[1]
port 924 nsew signal output
rlabel metal3 s 0 60800 800 60920 6 sb_hsize[2]
port 925 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 sb_htrans[0]
port 926 nsew signal output
rlabel metal3 s 0 61480 800 61600 6 sb_htrans[1]
port 927 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 sb_hwdata[0]
port 928 nsew signal output
rlabel metal3 s 0 65832 800 65952 6 sb_hwdata[10]
port 929 nsew signal output
rlabel metal3 s 0 66104 800 66224 6 sb_hwdata[11]
port 930 nsew signal output
rlabel metal3 s 0 66512 800 66632 6 sb_hwdata[12]
port 931 nsew signal output
rlabel metal3 s 0 66920 800 67040 6 sb_hwdata[13]
port 932 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 sb_hwdata[14]
port 933 nsew signal output
rlabel metal3 s 0 67600 800 67720 6 sb_hwdata[15]
port 934 nsew signal output
rlabel metal3 s 0 67872 800 67992 6 sb_hwdata[16]
port 935 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 sb_hwdata[17]
port 936 nsew signal output
rlabel metal3 s 0 68688 800 68808 6 sb_hwdata[18]
port 937 nsew signal output
rlabel metal3 s 0 68960 800 69080 6 sb_hwdata[19]
port 938 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 sb_hwdata[1]
port 939 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 sb_hwdata[20]
port 940 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 sb_hwdata[21]
port 941 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 sb_hwdata[22]
port 942 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 sb_hwdata[23]
port 943 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 sb_hwdata[24]
port 944 nsew signal output
rlabel metal3 s 0 71136 800 71256 6 sb_hwdata[25]
port 945 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 sb_hwdata[26]
port 946 nsew signal output
rlabel metal3 s 0 71816 800 71936 6 sb_hwdata[27]
port 947 nsew signal output
rlabel metal3 s 0 72224 800 72344 6 sb_hwdata[28]
port 948 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 sb_hwdata[29]
port 949 nsew signal output
rlabel metal3 s 0 62976 800 63096 6 sb_hwdata[2]
port 950 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 sb_hwdata[30]
port 951 nsew signal output
rlabel metal3 s 0 73312 800 73432 6 sb_hwdata[31]
port 952 nsew signal output
rlabel metal3 s 0 73584 800 73704 6 sb_hwdata[32]
port 953 nsew signal output
rlabel metal3 s 0 73992 800 74112 6 sb_hwdata[33]
port 954 nsew signal output
rlabel metal3 s 0 74400 800 74520 6 sb_hwdata[34]
port 955 nsew signal output
rlabel metal3 s 0 74672 800 74792 6 sb_hwdata[35]
port 956 nsew signal output
rlabel metal3 s 0 75080 800 75200 6 sb_hwdata[36]
port 957 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 sb_hwdata[37]
port 958 nsew signal output
rlabel metal3 s 0 75760 800 75880 6 sb_hwdata[38]
port 959 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 sb_hwdata[39]
port 960 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 sb_hwdata[3]
port 961 nsew signal output
rlabel metal3 s 0 76576 800 76696 6 sb_hwdata[40]
port 962 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 sb_hwdata[41]
port 963 nsew signal output
rlabel metal3 s 0 77256 800 77376 6 sb_hwdata[42]
port 964 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 sb_hwdata[43]
port 965 nsew signal output
rlabel metal3 s 0 77936 800 78056 6 sb_hwdata[44]
port 966 nsew signal output
rlabel metal3 s 0 78344 800 78464 6 sb_hwdata[45]
port 967 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 sb_hwdata[46]
port 968 nsew signal output
rlabel metal3 s 0 79024 800 79144 6 sb_hwdata[47]
port 969 nsew signal output
rlabel metal3 s 0 79432 800 79552 6 sb_hwdata[48]
port 970 nsew signal output
rlabel metal3 s 0 79704 800 79824 6 sb_hwdata[49]
port 971 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 sb_hwdata[4]
port 972 nsew signal output
rlabel metal3 s 0 80112 800 80232 6 sb_hwdata[50]
port 973 nsew signal output
rlabel metal3 s 0 80384 800 80504 6 sb_hwdata[51]
port 974 nsew signal output
rlabel metal3 s 0 80792 800 80912 6 sb_hwdata[52]
port 975 nsew signal output
rlabel metal3 s 0 81200 800 81320 6 sb_hwdata[53]
port 976 nsew signal output
rlabel metal3 s 0 81472 800 81592 6 sb_hwdata[54]
port 977 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 sb_hwdata[55]
port 978 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 sb_hwdata[56]
port 979 nsew signal output
rlabel metal3 s 0 82560 800 82680 6 sb_hwdata[57]
port 980 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 sb_hwdata[58]
port 981 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 sb_hwdata[59]
port 982 nsew signal output
rlabel metal3 s 0 64064 800 64184 6 sb_hwdata[5]
port 983 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 sb_hwdata[60]
port 984 nsew signal output
rlabel metal3 s 0 84056 800 84176 6 sb_hwdata[61]
port 985 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 sb_hwdata[62]
port 986 nsew signal output
rlabel metal3 s 0 84736 800 84856 6 sb_hwdata[63]
port 987 nsew signal output
rlabel metal3 s 0 64336 800 64456 6 sb_hwdata[6]
port 988 nsew signal output
rlabel metal3 s 0 64744 800 64864 6 sb_hwdata[7]
port 989 nsew signal output
rlabel metal3 s 0 65016 800 65136 6 sb_hwdata[8]
port 990 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 sb_hwdata[9]
port 991 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 sb_hwrite
port 992 nsew signal output
rlabel metal3 s 0 262216 800 262336 6 scan_mode
port 993 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 soft_int
port 994 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 timer_int
port 995 nsew signal input
rlabel metal3 s 0 262896 800 263016 6 trace_rv_i_address_ip[0]
port 996 nsew signal output
rlabel metal3 s 0 266568 800 266688 6 trace_rv_i_address_ip[10]
port 997 nsew signal output
rlabel metal3 s 0 266840 800 266960 6 trace_rv_i_address_ip[11]
port 998 nsew signal output
rlabel metal3 s 0 267248 800 267368 6 trace_rv_i_address_ip[12]
port 999 nsew signal output
rlabel metal3 s 0 267656 800 267776 6 trace_rv_i_address_ip[13]
port 1000 nsew signal output
rlabel metal3 s 0 267928 800 268048 6 trace_rv_i_address_ip[14]
port 1001 nsew signal output
rlabel metal3 s 0 268336 800 268456 6 trace_rv_i_address_ip[15]
port 1002 nsew signal output
rlabel metal3 s 0 268608 800 268728 6 trace_rv_i_address_ip[16]
port 1003 nsew signal output
rlabel metal3 s 0 269016 800 269136 6 trace_rv_i_address_ip[17]
port 1004 nsew signal output
rlabel metal3 s 0 269424 800 269544 6 trace_rv_i_address_ip[18]
port 1005 nsew signal output
rlabel metal3 s 0 269696 800 269816 6 trace_rv_i_address_ip[19]
port 1006 nsew signal output
rlabel metal3 s 0 263304 800 263424 6 trace_rv_i_address_ip[1]
port 1007 nsew signal output
rlabel metal3 s 0 270104 800 270224 6 trace_rv_i_address_ip[20]
port 1008 nsew signal output
rlabel metal3 s 0 270512 800 270632 6 trace_rv_i_address_ip[21]
port 1009 nsew signal output
rlabel metal3 s 0 270784 800 270904 6 trace_rv_i_address_ip[22]
port 1010 nsew signal output
rlabel metal3 s 0 271192 800 271312 6 trace_rv_i_address_ip[23]
port 1011 nsew signal output
rlabel metal3 s 0 271464 800 271584 6 trace_rv_i_address_ip[24]
port 1012 nsew signal output
rlabel metal3 s 0 271872 800 271992 6 trace_rv_i_address_ip[25]
port 1013 nsew signal output
rlabel metal3 s 0 272280 800 272400 6 trace_rv_i_address_ip[26]
port 1014 nsew signal output
rlabel metal3 s 0 272552 800 272672 6 trace_rv_i_address_ip[27]
port 1015 nsew signal output
rlabel metal3 s 0 272960 800 273080 6 trace_rv_i_address_ip[28]
port 1016 nsew signal output
rlabel metal3 s 0 273368 800 273488 6 trace_rv_i_address_ip[29]
port 1017 nsew signal output
rlabel metal3 s 0 263712 800 263832 6 trace_rv_i_address_ip[2]
port 1018 nsew signal output
rlabel metal3 s 0 273640 800 273760 6 trace_rv_i_address_ip[30]
port 1019 nsew signal output
rlabel metal3 s 0 274048 800 274168 6 trace_rv_i_address_ip[31]
port 1020 nsew signal output
rlabel metal3 s 0 263984 800 264104 6 trace_rv_i_address_ip[3]
port 1021 nsew signal output
rlabel metal3 s 0 264392 800 264512 6 trace_rv_i_address_ip[4]
port 1022 nsew signal output
rlabel metal3 s 0 264800 800 264920 6 trace_rv_i_address_ip[5]
port 1023 nsew signal output
rlabel metal3 s 0 265072 800 265192 6 trace_rv_i_address_ip[6]
port 1024 nsew signal output
rlabel metal3 s 0 265480 800 265600 6 trace_rv_i_address_ip[7]
port 1025 nsew signal output
rlabel metal3 s 0 265752 800 265872 6 trace_rv_i_address_ip[8]
port 1026 nsew signal output
rlabel metal3 s 0 266160 800 266280 6 trace_rv_i_address_ip[9]
port 1027 nsew signal output
rlabel metal3 s 0 274320 800 274440 6 trace_rv_i_ecause_ip[0]
port 1028 nsew signal output
rlabel metal3 s 0 274728 800 274848 6 trace_rv_i_ecause_ip[1]
port 1029 nsew signal output
rlabel metal3 s 0 275136 800 275256 6 trace_rv_i_ecause_ip[2]
port 1030 nsew signal output
rlabel metal3 s 0 275408 800 275528 6 trace_rv_i_ecause_ip[3]
port 1031 nsew signal output
rlabel metal3 s 0 275816 800 275936 6 trace_rv_i_ecause_ip[4]
port 1032 nsew signal output
rlabel metal3 s 0 276224 800 276344 6 trace_rv_i_exception_ip
port 1033 nsew signal output
rlabel metal3 s 0 276496 800 276616 6 trace_rv_i_insn_ip[0]
port 1034 nsew signal output
rlabel metal3 s 0 280032 800 280152 6 trace_rv_i_insn_ip[10]
port 1035 nsew signal output
rlabel metal3 s 0 280440 800 280560 6 trace_rv_i_insn_ip[11]
port 1036 nsew signal output
rlabel metal3 s 0 280848 800 280968 6 trace_rv_i_insn_ip[12]
port 1037 nsew signal output
rlabel metal3 s 0 281120 800 281240 6 trace_rv_i_insn_ip[13]
port 1038 nsew signal output
rlabel metal3 s 0 281528 800 281648 6 trace_rv_i_insn_ip[14]
port 1039 nsew signal output
rlabel metal3 s 0 281936 800 282056 6 trace_rv_i_insn_ip[15]
port 1040 nsew signal output
rlabel metal3 s 0 282208 800 282328 6 trace_rv_i_insn_ip[16]
port 1041 nsew signal output
rlabel metal3 s 0 282616 800 282736 6 trace_rv_i_insn_ip[17]
port 1042 nsew signal output
rlabel metal3 s 0 282888 800 283008 6 trace_rv_i_insn_ip[18]
port 1043 nsew signal output
rlabel metal3 s 0 283296 800 283416 6 trace_rv_i_insn_ip[19]
port 1044 nsew signal output
rlabel metal3 s 0 276904 800 277024 6 trace_rv_i_insn_ip[1]
port 1045 nsew signal output
rlabel metal3 s 0 283704 800 283824 6 trace_rv_i_insn_ip[20]
port 1046 nsew signal output
rlabel metal3 s 0 283976 800 284096 6 trace_rv_i_insn_ip[21]
port 1047 nsew signal output
rlabel metal3 s 0 284384 800 284504 6 trace_rv_i_insn_ip[22]
port 1048 nsew signal output
rlabel metal3 s 0 284792 800 284912 6 trace_rv_i_insn_ip[23]
port 1049 nsew signal output
rlabel metal3 s 0 285064 800 285184 6 trace_rv_i_insn_ip[24]
port 1050 nsew signal output
rlabel metal3 s 0 285472 800 285592 6 trace_rv_i_insn_ip[25]
port 1051 nsew signal output
rlabel metal3 s 0 285744 800 285864 6 trace_rv_i_insn_ip[26]
port 1052 nsew signal output
rlabel metal3 s 0 286152 800 286272 6 trace_rv_i_insn_ip[27]
port 1053 nsew signal output
rlabel metal3 s 0 286560 800 286680 6 trace_rv_i_insn_ip[28]
port 1054 nsew signal output
rlabel metal3 s 0 286832 800 286952 6 trace_rv_i_insn_ip[29]
port 1055 nsew signal output
rlabel metal3 s 0 277176 800 277296 6 trace_rv_i_insn_ip[2]
port 1056 nsew signal output
rlabel metal3 s 0 287240 800 287360 6 trace_rv_i_insn_ip[30]
port 1057 nsew signal output
rlabel metal3 s 0 287648 800 287768 6 trace_rv_i_insn_ip[31]
port 1058 nsew signal output
rlabel metal3 s 0 277584 800 277704 6 trace_rv_i_insn_ip[3]
port 1059 nsew signal output
rlabel metal3 s 0 277992 800 278112 6 trace_rv_i_insn_ip[4]
port 1060 nsew signal output
rlabel metal3 s 0 278264 800 278384 6 trace_rv_i_insn_ip[5]
port 1061 nsew signal output
rlabel metal3 s 0 278672 800 278792 6 trace_rv_i_insn_ip[6]
port 1062 nsew signal output
rlabel metal3 s 0 279080 800 279200 6 trace_rv_i_insn_ip[7]
port 1063 nsew signal output
rlabel metal3 s 0 279352 800 279472 6 trace_rv_i_insn_ip[8]
port 1064 nsew signal output
rlabel metal3 s 0 279760 800 279880 6 trace_rv_i_insn_ip[9]
port 1065 nsew signal output
rlabel metal3 s 0 287920 800 288040 6 trace_rv_i_interrupt_ip
port 1066 nsew signal output
rlabel metal3 s 0 288328 800 288448 6 trace_rv_i_tval_ip[0]
port 1067 nsew signal output
rlabel metal3 s 0 291864 800 291984 6 trace_rv_i_tval_ip[10]
port 1068 nsew signal output
rlabel metal3 s 0 292272 800 292392 6 trace_rv_i_tval_ip[11]
port 1069 nsew signal output
rlabel metal3 s 0 292544 800 292664 6 trace_rv_i_tval_ip[12]
port 1070 nsew signal output
rlabel metal3 s 0 292952 800 293072 6 trace_rv_i_tval_ip[13]
port 1071 nsew signal output
rlabel metal3 s 0 293360 800 293480 6 trace_rv_i_tval_ip[14]
port 1072 nsew signal output
rlabel metal3 s 0 293632 800 293752 6 trace_rv_i_tval_ip[15]
port 1073 nsew signal output
rlabel metal3 s 0 294040 800 294160 6 trace_rv_i_tval_ip[16]
port 1074 nsew signal output
rlabel metal3 s 0 294312 800 294432 6 trace_rv_i_tval_ip[17]
port 1075 nsew signal output
rlabel metal3 s 0 294720 800 294840 6 trace_rv_i_tval_ip[18]
port 1076 nsew signal output
rlabel metal3 s 0 295128 800 295248 6 trace_rv_i_tval_ip[19]
port 1077 nsew signal output
rlabel metal3 s 0 288600 800 288720 6 trace_rv_i_tval_ip[1]
port 1078 nsew signal output
rlabel metal3 s 0 295400 800 295520 6 trace_rv_i_tval_ip[20]
port 1079 nsew signal output
rlabel metal3 s 0 295808 800 295928 6 trace_rv_i_tval_ip[21]
port 1080 nsew signal output
rlabel metal3 s 0 296216 800 296336 6 trace_rv_i_tval_ip[22]
port 1081 nsew signal output
rlabel metal3 s 0 296488 800 296608 6 trace_rv_i_tval_ip[23]
port 1082 nsew signal output
rlabel metal3 s 0 296896 800 297016 6 trace_rv_i_tval_ip[24]
port 1083 nsew signal output
rlabel metal3 s 0 297168 800 297288 6 trace_rv_i_tval_ip[25]
port 1084 nsew signal output
rlabel metal3 s 0 297576 800 297696 6 trace_rv_i_tval_ip[26]
port 1085 nsew signal output
rlabel metal3 s 0 297984 800 298104 6 trace_rv_i_tval_ip[27]
port 1086 nsew signal output
rlabel metal3 s 0 298256 800 298376 6 trace_rv_i_tval_ip[28]
port 1087 nsew signal output
rlabel metal3 s 0 298664 800 298784 6 trace_rv_i_tval_ip[29]
port 1088 nsew signal output
rlabel metal3 s 0 289008 800 289128 6 trace_rv_i_tval_ip[2]
port 1089 nsew signal output
rlabel metal3 s 0 299072 800 299192 6 trace_rv_i_tval_ip[30]
port 1090 nsew signal output
rlabel metal3 s 0 299344 800 299464 6 trace_rv_i_tval_ip[31]
port 1091 nsew signal output
rlabel metal3 s 0 289416 800 289536 6 trace_rv_i_tval_ip[3]
port 1092 nsew signal output
rlabel metal3 s 0 289688 800 289808 6 trace_rv_i_tval_ip[4]
port 1093 nsew signal output
rlabel metal3 s 0 290096 800 290216 6 trace_rv_i_tval_ip[5]
port 1094 nsew signal output
rlabel metal3 s 0 290504 800 290624 6 trace_rv_i_tval_ip[6]
port 1095 nsew signal output
rlabel metal3 s 0 290776 800 290896 6 trace_rv_i_tval_ip[7]
port 1096 nsew signal output
rlabel metal3 s 0 291184 800 291304 6 trace_rv_i_tval_ip[8]
port 1097 nsew signal output
rlabel metal3 s 0 291456 800 291576 6 trace_rv_i_tval_ip[9]
port 1098 nsew signal output
rlabel metal3 s 0 299752 800 299872 6 trace_rv_i_valid_ip
port 1099 nsew signal output
rlabel metal4 s 249968 2128 250288 297616 6 VPWR
port 1100 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 297616 6 VPWR
port 1101 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 297616 6 VPWR
port 1102 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 297616 6 VPWR
port 1103 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 297616 6 VPWR
port 1104 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 297616 6 VPWR
port 1105 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 297616 6 VPWR
port 1106 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 297616 6 VPWR
port 1107 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 297616 6 VPWR
port 1108 nsew power bidirectional
rlabel metal4 s 265328 2128 265648 297616 6 VGND
port 1109 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 297616 6 VGND
port 1110 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 297616 6 VGND
port 1111 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 297616 6 VGND
port 1112 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 297616 6 VGND
port 1113 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 297616 6 VGND
port 1114 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 297616 6 VGND
port 1115 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 297616 6 VGND
port 1116 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 297616 6 VGND
port 1117 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 279390 299872
string LEFview TRUE
<< end >>
