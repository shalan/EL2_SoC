VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM_4K
  CLASS BLOCK ;
  FOREIGN DFFRAM_4K ;
  ORIGIN 0.000 0.000 ;
  SIZE 1159.120 BY 1489.360 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.480 1485.360 469.760 1489.360 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.740 1485.360 484.020 1489.360 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.460 1485.360 498.740 1489.360 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.180 1485.360 513.460 1489.360 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.900 1485.360 528.180 1489.360 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.620 1485.360 542.900 1489.360 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.880 1485.360 557.160 1489.360 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.600 1485.360 571.880 1489.360 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.320 1485.360 586.600 1489.360 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.040 1485.360 601.320 1489.360 ;
    END
  END A[9]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.760 1485.360 616.040 1489.360 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.160 1485.360 703.440 1489.360 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.440 1485.360 849.720 1489.360 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.160 1485.360 864.440 1489.360 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.880 1485.360 879.160 1489.360 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.600 1485.360 893.880 1489.360 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.860 1485.360 908.140 1489.360 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.580 1485.360 922.860 1489.360 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.300 1485.360 937.580 1489.360 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.020 1485.360 952.300 1489.360 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.280 1485.360 966.560 1489.360 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.000 1485.360 981.280 1489.360 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.880 1485.360 718.160 1489.360 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.720 1485.360 996.000 1489.360 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.440 1485.360 1010.720 1489.360 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.160 1485.360 1025.440 1489.360 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.420 1485.360 1039.700 1489.360 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.140 1485.360 1054.420 1489.360 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.860 1485.360 1069.140 1489.360 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.580 1485.360 1083.860 1489.360 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.300 1485.360 1098.580 1489.360 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.560 1485.360 1112.840 1489.360 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.280 1485.360 1127.560 1489.360 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.600 1485.360 732.880 1489.360 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.000 1485.360 1142.280 1489.360 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.720 1485.360 1157.000 1489.360 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.320 1485.360 747.600 1489.360 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.580 1485.360 761.860 1489.360 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.300 1485.360 776.580 1489.360 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.020 1485.360 791.300 1489.360 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.740 1485.360 806.020 1489.360 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.460 1485.360 820.740 1489.360 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.720 1485.360 835.000 1489.360 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.660 1485.360 1.940 1489.360 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.480 1485.360 147.760 1489.360 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.200 1485.360 162.480 1489.360 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.920 1485.360 177.200 1489.360 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.640 1485.360 191.920 1489.360 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.360 1485.360 206.640 1489.360 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.620 1485.360 220.900 1489.360 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.340 1485.360 235.620 1489.360 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.060 1485.360 250.340 1489.360 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.780 1485.360 265.060 1489.360 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.040 1485.360 279.320 1489.360 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.920 1485.360 16.200 1489.360 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.760 1485.360 294.040 1489.360 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.480 1485.360 308.760 1489.360 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.200 1485.360 323.480 1489.360 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.920 1485.360 338.200 1489.360 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.180 1485.360 352.460 1489.360 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.900 1485.360 367.180 1489.360 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.620 1485.360 381.900 1489.360 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.340 1485.360 396.620 1489.360 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.060 1485.360 411.340 1489.360 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.320 1485.360 425.600 1489.360 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.640 1485.360 30.920 1489.360 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.040 1485.360 440.320 1489.360 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.760 1485.360 455.040 1489.360 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.360 1485.360 45.640 1489.360 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.080 1485.360 60.360 1489.360 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.340 1485.360 74.620 1489.360 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.060 1485.360 89.340 1489.360 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.780 1485.360 104.060 1489.360 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.500 1485.360 118.780 1489.360 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.220 1485.360 133.500 1489.360 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.900 1485.360 689.180 1489.360 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.020 1485.360 630.300 1489.360 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.740 1485.360 645.020 1489.360 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.460 1485.360 659.740 1489.360 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.180 1485.360 674.460 1489.360 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1095.710 0.000 1097.310 1477.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 975.710 0.000 977.310 1477.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 855.710 0.000 857.310 1477.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 735.710 0.000 737.310 1477.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 615.710 0.000 617.310 1477.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 495.710 0.000 497.310 1477.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 375.710 0.000 377.310 1477.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 255.710 0.000 257.310 1477.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 135.710 0.000 137.310 1477.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.710 0.000 17.310 1477.440 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1155.710 0.000 1157.310 1477.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1035.710 0.000 1037.310 1477.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 915.710 0.000 917.310 1477.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 795.710 0.000 797.310 1477.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 675.710 0.000 677.310 1477.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 555.710 0.000 557.310 1477.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 435.710 0.000 437.310 1477.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 315.710 0.000 317.310 1477.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 195.710 0.000 197.310 1477.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 75.710 0.000 77.310 1477.440 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.190 0.155 1158.930 1477.285 ;
      LAYER met1 ;
        RECT 0.190 0.000 1158.930 1478.860 ;
      LAYER met2 ;
        RECT 2.220 1485.080 15.640 1485.360 ;
        RECT 16.480 1485.080 30.360 1485.360 ;
        RECT 31.200 1485.080 45.080 1485.360 ;
        RECT 45.920 1485.080 59.800 1485.360 ;
        RECT 60.640 1485.080 74.060 1485.360 ;
        RECT 74.900 1485.080 88.780 1485.360 ;
        RECT 89.620 1485.080 103.500 1485.360 ;
        RECT 104.340 1485.080 118.220 1485.360 ;
        RECT 119.060 1485.080 132.940 1485.360 ;
        RECT 133.780 1485.080 147.200 1485.360 ;
        RECT 148.040 1485.080 161.920 1485.360 ;
        RECT 162.760 1485.080 176.640 1485.360 ;
        RECT 177.480 1485.080 191.360 1485.360 ;
        RECT 192.200 1485.080 206.080 1485.360 ;
        RECT 206.920 1485.080 220.340 1485.360 ;
        RECT 221.180 1485.080 235.060 1485.360 ;
        RECT 235.900 1485.080 249.780 1485.360 ;
        RECT 250.620 1485.080 264.500 1485.360 ;
        RECT 265.340 1485.080 278.760 1485.360 ;
        RECT 279.600 1485.080 293.480 1485.360 ;
        RECT 294.320 1485.080 308.200 1485.360 ;
        RECT 309.040 1485.080 322.920 1485.360 ;
        RECT 323.760 1485.080 337.640 1485.360 ;
        RECT 338.480 1485.080 351.900 1485.360 ;
        RECT 352.740 1485.080 366.620 1485.360 ;
        RECT 367.460 1485.080 381.340 1485.360 ;
        RECT 382.180 1485.080 396.060 1485.360 ;
        RECT 396.900 1485.080 410.780 1485.360 ;
        RECT 411.620 1485.080 425.040 1485.360 ;
        RECT 425.880 1485.080 439.760 1485.360 ;
        RECT 440.600 1485.080 454.480 1485.360 ;
        RECT 455.320 1485.080 469.200 1485.360 ;
        RECT 470.040 1485.080 483.460 1485.360 ;
        RECT 484.300 1485.080 498.180 1485.360 ;
        RECT 499.020 1485.080 512.900 1485.360 ;
        RECT 513.740 1485.080 527.620 1485.360 ;
        RECT 528.460 1485.080 542.340 1485.360 ;
        RECT 543.180 1485.080 556.600 1485.360 ;
        RECT 557.440 1485.080 571.320 1485.360 ;
        RECT 572.160 1485.080 586.040 1485.360 ;
        RECT 586.880 1485.080 600.760 1485.360 ;
        RECT 601.600 1485.080 615.480 1485.360 ;
        RECT 616.320 1485.080 629.740 1485.360 ;
        RECT 630.580 1485.080 644.460 1485.360 ;
        RECT 645.300 1485.080 659.180 1485.360 ;
        RECT 660.020 1485.080 673.900 1485.360 ;
        RECT 674.740 1485.080 688.620 1485.360 ;
        RECT 689.460 1485.080 702.880 1485.360 ;
        RECT 703.720 1485.080 717.600 1485.360 ;
        RECT 718.440 1485.080 732.320 1485.360 ;
        RECT 733.160 1485.080 747.040 1485.360 ;
        RECT 747.880 1485.080 761.300 1485.360 ;
        RECT 762.140 1485.080 776.020 1485.360 ;
        RECT 776.860 1485.080 790.740 1485.360 ;
        RECT 791.580 1485.080 805.460 1485.360 ;
        RECT 806.300 1485.080 820.180 1485.360 ;
        RECT 821.020 1485.080 834.440 1485.360 ;
        RECT 835.280 1485.080 849.160 1485.360 ;
        RECT 850.000 1485.080 863.880 1485.360 ;
        RECT 864.720 1485.080 878.600 1485.360 ;
        RECT 879.440 1485.080 893.320 1485.360 ;
        RECT 894.160 1485.080 907.580 1485.360 ;
        RECT 908.420 1485.080 922.300 1485.360 ;
        RECT 923.140 1485.080 937.020 1485.360 ;
        RECT 937.860 1485.080 951.740 1485.360 ;
        RECT 952.580 1485.080 966.000 1485.360 ;
        RECT 966.840 1485.080 980.720 1485.360 ;
        RECT 981.560 1485.080 995.440 1485.360 ;
        RECT 996.280 1485.080 1010.160 1485.360 ;
        RECT 1011.000 1485.080 1024.880 1485.360 ;
        RECT 1025.720 1485.080 1039.140 1485.360 ;
        RECT 1039.980 1485.080 1053.860 1485.360 ;
        RECT 1054.700 1485.080 1068.580 1485.360 ;
        RECT 1069.420 1485.080 1083.300 1485.360 ;
        RECT 1084.140 1485.080 1098.020 1485.360 ;
        RECT 1098.860 1485.080 1112.280 1485.360 ;
        RECT 1113.120 1485.080 1127.000 1485.360 ;
        RECT 1127.840 1485.080 1141.720 1485.360 ;
        RECT 1142.560 1485.080 1156.440 1485.360 ;
        RECT 1157.280 1485.080 1157.910 1485.360 ;
        RECT 1.670 0.000 1157.910 1485.080 ;
      LAYER met3 ;
        RECT 3.015 0.075 1157.310 1477.365 ;
      LAYER met4 ;
        RECT 20.725 42.575 75.310 1474.985 ;
        RECT 77.710 42.575 135.310 1474.985 ;
        RECT 137.710 42.575 195.310 1474.985 ;
        RECT 197.710 42.575 255.310 1474.985 ;
        RECT 257.710 42.575 315.310 1474.985 ;
        RECT 317.710 42.575 375.310 1474.985 ;
        RECT 377.710 42.575 435.310 1474.985 ;
        RECT 437.710 42.575 495.310 1474.985 ;
        RECT 497.710 42.575 555.310 1474.985 ;
        RECT 557.710 42.575 615.310 1474.985 ;
        RECT 617.710 42.575 675.310 1474.985 ;
        RECT 677.710 42.575 735.310 1474.985 ;
        RECT 737.710 42.575 795.310 1474.985 ;
        RECT 797.710 42.575 855.310 1474.985 ;
        RECT 857.710 42.575 915.310 1474.985 ;
        RECT 917.710 42.575 975.310 1474.985 ;
        RECT 977.710 42.575 1035.310 1474.985 ;
        RECT 1037.710 42.575 1095.310 1474.985 ;
        RECT 1097.710 42.575 1140.695 1474.985 ;
        RECT 15.710 0.300 1157.310 1477.440 ;
  END
END DFFRAM_4K
END LIBRARY

