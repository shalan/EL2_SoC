VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO el2_swerv_wrapper
  CLASS BLOCK ;
  FOREIGN el2_swerv_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 1396.950 BY 1499.360 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END clk
  PIN core_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1239.680 4.000 1240.280 ;
    END
  END core_id[0]
  PIN core_id[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1257.360 4.000 1257.960 ;
    END
  END core_id[10]
  PIN core_id[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1259.400 4.000 1260.000 ;
    END
  END core_id[11]
  PIN core_id[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1261.440 4.000 1262.040 ;
    END
  END core_id[12]
  PIN core_id[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1262.800 4.000 1263.400 ;
    END
  END core_id[13]
  PIN core_id[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.840 4.000 1265.440 ;
    END
  END core_id[14]
  PIN core_id[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1266.200 4.000 1266.800 ;
    END
  END core_id[15]
  PIN core_id[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.240 4.000 1268.840 ;
    END
  END core_id[16]
  PIN core_id[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1270.280 4.000 1270.880 ;
    END
  END core_id[17]
  PIN core_id[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1271.640 4.000 1272.240 ;
    END
  END core_id[18]
  PIN core_id[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1273.680 4.000 1274.280 ;
    END
  END core_id[19]
  PIN core_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.720 4.000 1242.320 ;
    END
  END core_id[1]
  PIN core_id[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.720 4.000 1276.320 ;
    END
  END core_id[20]
  PIN core_id[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1277.080 4.000 1277.680 ;
    END
  END core_id[21]
  PIN core_id[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1279.120 4.000 1279.720 ;
    END
  END core_id[22]
  PIN core_id[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1280.480 4.000 1281.080 ;
    END
  END core_id[23]
  PIN core_id[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1282.520 4.000 1283.120 ;
    END
  END core_id[24]
  PIN core_id[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1284.560 4.000 1285.160 ;
    END
  END core_id[25]
  PIN core_id[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.920 4.000 1286.520 ;
    END
  END core_id[26]
  PIN core_id[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1287.960 4.000 1288.560 ;
    END
  END core_id[27]
  PIN core_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.080 4.000 1243.680 ;
    END
  END core_id[2]
  PIN core_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1245.120 4.000 1245.720 ;
    END
  END core_id[3]
  PIN core_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.160 4.000 1247.760 ;
    END
  END core_id[4]
  PIN core_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1248.520 4.000 1249.120 ;
    END
  END core_id[5]
  PIN core_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1250.560 4.000 1251.160 ;
    END
  END core_id[6]
  PIN core_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1251.920 4.000 1252.520 ;
    END
  END core_id[7]
  PIN core_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1253.960 4.000 1254.560 ;
    END
  END core_id[8]
  PIN core_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1256.000 4.000 1256.600 ;
    END
  END core_id[9]
  PIN dbg_bus_clk_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END dbg_bus_clk_en
  PIN dbg_rst_l
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END dbg_rst_l
  PIN dccm_ext_in_pkt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 868.400 4.000 869.000 ;
    END
  END dccm_ext_in_pkt[0]
  PIN dccm_ext_in_pkt[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.080 4.000 886.680 ;
    END
  END dccm_ext_in_pkt[10]
  PIN dccm_ext_in_pkt[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END dccm_ext_in_pkt[11]
  PIN dccm_ext_in_pkt[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 889.480 4.000 890.080 ;
    END
  END dccm_ext_in_pkt[12]
  PIN dccm_ext_in_pkt[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 891.520 4.000 892.120 ;
    END
  END dccm_ext_in_pkt[13]
  PIN dccm_ext_in_pkt[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END dccm_ext_in_pkt[14]
  PIN dccm_ext_in_pkt[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.920 4.000 895.520 ;
    END
  END dccm_ext_in_pkt[15]
  PIN dccm_ext_in_pkt[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.960 4.000 897.560 ;
    END
  END dccm_ext_in_pkt[16]
  PIN dccm_ext_in_pkt[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 898.320 4.000 898.920 ;
    END
  END dccm_ext_in_pkt[17]
  PIN dccm_ext_in_pkt[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 900.360 4.000 900.960 ;
    END
  END dccm_ext_in_pkt[18]
  PIN dccm_ext_in_pkt[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 902.400 4.000 903.000 ;
    END
  END dccm_ext_in_pkt[19]
  PIN dccm_ext_in_pkt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 869.760 4.000 870.360 ;
    END
  END dccm_ext_in_pkt[1]
  PIN dccm_ext_in_pkt[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.760 4.000 904.360 ;
    END
  END dccm_ext_in_pkt[20]
  PIN dccm_ext_in_pkt[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END dccm_ext_in_pkt[21]
  PIN dccm_ext_in_pkt[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END dccm_ext_in_pkt[22]
  PIN dccm_ext_in_pkt[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.200 4.000 909.800 ;
    END
  END dccm_ext_in_pkt[23]
  PIN dccm_ext_in_pkt[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END dccm_ext_in_pkt[24]
  PIN dccm_ext_in_pkt[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 912.600 4.000 913.200 ;
    END
  END dccm_ext_in_pkt[25]
  PIN dccm_ext_in_pkt[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END dccm_ext_in_pkt[26]
  PIN dccm_ext_in_pkt[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.680 4.000 917.280 ;
    END
  END dccm_ext_in_pkt[27]
  PIN dccm_ext_in_pkt[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END dccm_ext_in_pkt[28]
  PIN dccm_ext_in_pkt[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.080 4.000 920.680 ;
    END
  END dccm_ext_in_pkt[29]
  PIN dccm_ext_in_pkt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.800 4.000 872.400 ;
    END
  END dccm_ext_in_pkt[2]
  PIN dccm_ext_in_pkt[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 922.120 4.000 922.720 ;
    END
  END dccm_ext_in_pkt[30]
  PIN dccm_ext_in_pkt[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 923.480 4.000 924.080 ;
    END
  END dccm_ext_in_pkt[31]
  PIN dccm_ext_in_pkt[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 925.520 4.000 926.120 ;
    END
  END dccm_ext_in_pkt[32]
  PIN dccm_ext_in_pkt[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.880 4.000 927.480 ;
    END
  END dccm_ext_in_pkt[33]
  PIN dccm_ext_in_pkt[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.920 4.000 929.520 ;
    END
  END dccm_ext_in_pkt[34]
  PIN dccm_ext_in_pkt[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END dccm_ext_in_pkt[35]
  PIN dccm_ext_in_pkt[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 932.320 4.000 932.920 ;
    END
  END dccm_ext_in_pkt[36]
  PIN dccm_ext_in_pkt[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 934.360 4.000 934.960 ;
    END
  END dccm_ext_in_pkt[37]
  PIN dccm_ext_in_pkt[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 936.400 4.000 937.000 ;
    END
  END dccm_ext_in_pkt[38]
  PIN dccm_ext_in_pkt[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.760 4.000 938.360 ;
    END
  END dccm_ext_in_pkt[39]
  PIN dccm_ext_in_pkt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END dccm_ext_in_pkt[3]
  PIN dccm_ext_in_pkt[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.800 4.000 940.400 ;
    END
  END dccm_ext_in_pkt[40]
  PIN dccm_ext_in_pkt[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END dccm_ext_in_pkt[41]
  PIN dccm_ext_in_pkt[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.200 4.000 943.800 ;
    END
  END dccm_ext_in_pkt[42]
  PIN dccm_ext_in_pkt[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END dccm_ext_in_pkt[43]
  PIN dccm_ext_in_pkt[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 946.600 4.000 947.200 ;
    END
  END dccm_ext_in_pkt[44]
  PIN dccm_ext_in_pkt[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END dccm_ext_in_pkt[45]
  PIN dccm_ext_in_pkt[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.680 4.000 951.280 ;
    END
  END dccm_ext_in_pkt[46]
  PIN dccm_ext_in_pkt[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END dccm_ext_in_pkt[47]
  PIN dccm_ext_in_pkt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.200 4.000 875.800 ;
    END
  END dccm_ext_in_pkt[4]
  PIN dccm_ext_in_pkt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END dccm_ext_in_pkt[5]
  PIN dccm_ext_in_pkt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.280 4.000 879.880 ;
    END
  END dccm_ext_in_pkt[6]
  PIN dccm_ext_in_pkt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END dccm_ext_in_pkt[7]
  PIN dccm_ext_in_pkt[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 882.680 4.000 883.280 ;
    END
  END dccm_ext_in_pkt[8]
  PIN dccm_ext_in_pkt[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END dccm_ext_in_pkt[9]
  PIN debug_brkpt_status
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1298.840 4.000 1299.440 ;
    END
  END debug_brkpt_status
  PIN dec_tlu_perfcnt0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1168.280 4.000 1168.880 ;
    END
  END dec_tlu_perfcnt0
  PIN dec_tlu_perfcnt1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1170.320 4.000 1170.920 ;
    END
  END dec_tlu_perfcnt1
  PIN dec_tlu_perfcnt2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1171.680 4.000 1172.280 ;
    END
  END dec_tlu_perfcnt2
  PIN dec_tlu_perfcnt3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.720 4.000 1174.320 ;
    END
  END dec_tlu_perfcnt3
  PIN dma_bus_clk_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END dma_bus_clk_en
  PIN dma_haddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.720 4.000 545.320 ;
    END
  END dma_haddr[0]
  PIN dma_haddr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END dma_haddr[10]
  PIN dma_haddr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END dma_haddr[11]
  PIN dma_haddr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 566.480 4.000 567.080 ;
    END
  END dma_haddr[12]
  PIN dma_haddr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END dma_haddr[13]
  PIN dma_haddr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END dma_haddr[14]
  PIN dma_haddr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.920 4.000 572.520 ;
    END
  END dma_haddr[15]
  PIN dma_haddr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END dma_haddr[16]
  PIN dma_haddr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END dma_haddr[17]
  PIN dma_haddr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 577.360 4.000 577.960 ;
    END
  END dma_haddr[18]
  PIN dma_haddr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END dma_haddr[19]
  PIN dma_haddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END dma_haddr[1]
  PIN dma_haddr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END dma_haddr[20]
  PIN dma_haddr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.800 4.000 583.400 ;
    END
  END dma_haddr[21]
  PIN dma_haddr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.160 4.000 584.760 ;
    END
  END dma_haddr[22]
  PIN dma_haddr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END dma_haddr[23]
  PIN dma_haddr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END dma_haddr[24]
  PIN dma_haddr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 589.600 4.000 590.200 ;
    END
  END dma_haddr[25]
  PIN dma_haddr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END dma_haddr[26]
  PIN dma_haddr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END dma_haddr[27]
  PIN dma_haddr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END dma_haddr[28]
  PIN dma_haddr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END dma_haddr[29]
  PIN dma_haddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 4.000 549.400 ;
    END
  END dma_haddr[2]
  PIN dma_haddr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END dma_haddr[30]
  PIN dma_haddr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 600.480 4.000 601.080 ;
    END
  END dma_haddr[31]
  PIN dma_haddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.160 4.000 550.760 ;
    END
  END dma_haddr[3]
  PIN dma_haddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END dma_haddr[4]
  PIN dma_haddr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END dma_haddr[5]
  PIN dma_haddr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END dma_haddr[6]
  PIN dma_haddr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END dma_haddr[7]
  PIN dma_haddr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END dma_haddr[8]
  PIN dma_haddr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END dma_haddr[9]
  PIN dma_hburst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END dma_hburst[0]
  PIN dma_hburst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.880 4.000 604.480 ;
    END
  END dma_hburst[1]
  PIN dma_hburst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.920 4.000 606.520 ;
    END
  END dma_hburst[2]
  PIN dma_hmastlock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.280 4.000 607.880 ;
    END
  END dma_hmastlock
  PIN dma_hprot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END dma_hprot[0]
  PIN dma_hprot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 611.360 4.000 611.960 ;
    END
  END dma_hprot[1]
  PIN dma_hprot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.720 4.000 613.320 ;
    END
  END dma_hprot[2]
  PIN dma_hprot[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END dma_hprot[3]
  PIN dma_hrdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END dma_hrdata[0]
  PIN dma_hrdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.960 4.000 761.560 ;
    END
  END dma_hrdata[10]
  PIN dma_hrdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END dma_hrdata[11]
  PIN dma_hrdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END dma_hrdata[12]
  PIN dma_hrdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 766.400 4.000 767.000 ;
    END
  END dma_hrdata[13]
  PIN dma_hrdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END dma_hrdata[14]
  PIN dma_hrdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END dma_hrdata[15]
  PIN dma_hrdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END dma_hrdata[16]
  PIN dma_hrdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.880 4.000 774.480 ;
    END
  END dma_hrdata[17]
  PIN dma_hrdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END dma_hrdata[18]
  PIN dma_hrdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.280 4.000 777.880 ;
    END
  END dma_hrdata[19]
  PIN dma_hrdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.320 4.000 745.920 ;
    END
  END dma_hrdata[1]
  PIN dma_hrdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END dma_hrdata[20]
  PIN dma_hrdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END dma_hrdata[21]
  PIN dma_hrdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.720 4.000 783.320 ;
    END
  END dma_hrdata[22]
  PIN dma_hrdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.080 4.000 784.680 ;
    END
  END dma_hrdata[23]
  PIN dma_hrdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END dma_hrdata[24]
  PIN dma_hrdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.160 4.000 788.760 ;
    END
  END dma_hrdata[25]
  PIN dma_hrdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 789.520 4.000 790.120 ;
    END
  END dma_hrdata[26]
  PIN dma_hrdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 791.560 4.000 792.160 ;
    END
  END dma_hrdata[27]
  PIN dma_hrdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 793.600 4.000 794.200 ;
    END
  END dma_hrdata[28]
  PIN dma_hrdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.960 4.000 795.560 ;
    END
  END dma_hrdata[29]
  PIN dma_hrdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END dma_hrdata[2]
  PIN dma_hrdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END dma_hrdata[30]
  PIN dma_hrdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 798.360 4.000 798.960 ;
    END
  END dma_hrdata[31]
  PIN dma_hrdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 800.400 4.000 801.000 ;
    END
  END dma_hrdata[32]
  PIN dma_hrdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END dma_hrdata[33]
  PIN dma_hrdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.800 4.000 804.400 ;
    END
  END dma_hrdata[34]
  PIN dma_hrdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END dma_hrdata[35]
  PIN dma_hrdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END dma_hrdata[36]
  PIN dma_hrdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END dma_hrdata[37]
  PIN dma_hrdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.280 4.000 811.880 ;
    END
  END dma_hrdata[38]
  PIN dma_hrdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END dma_hrdata[39]
  PIN dma_hrdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.720 4.000 749.320 ;
    END
  END dma_hrdata[3]
  PIN dma_hrdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END dma_hrdata[40]
  PIN dma_hrdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.720 4.000 817.320 ;
    END
  END dma_hrdata[41]
  PIN dma_hrdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.080 4.000 818.680 ;
    END
  END dma_hrdata[42]
  PIN dma_hrdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.120 4.000 820.720 ;
    END
  END dma_hrdata[43]
  PIN dma_hrdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.160 4.000 822.760 ;
    END
  END dma_hrdata[44]
  PIN dma_hrdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 823.520 4.000 824.120 ;
    END
  END dma_hrdata[45]
  PIN dma_hrdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END dma_hrdata[46]
  PIN dma_hrdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.920 4.000 827.520 ;
    END
  END dma_hrdata[47]
  PIN dma_hrdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.960 4.000 829.560 ;
    END
  END dma_hrdata[48]
  PIN dma_hrdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 831.000 4.000 831.600 ;
    END
  END dma_hrdata[49]
  PIN dma_hrdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.760 4.000 751.360 ;
    END
  END dma_hrdata[4]
  PIN dma_hrdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END dma_hrdata[50]
  PIN dma_hrdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 834.400 4.000 835.000 ;
    END
  END dma_hrdata[51]
  PIN dma_hrdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END dma_hrdata[52]
  PIN dma_hrdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END dma_hrdata[53]
  PIN dma_hrdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END dma_hrdata[54]
  PIN dma_hrdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 841.200 4.000 841.800 ;
    END
  END dma_hrdata[55]
  PIN dma_hrdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END dma_hrdata[56]
  PIN dma_hrdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.280 4.000 845.880 ;
    END
  END dma_hrdata[57]
  PIN dma_hrdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END dma_hrdata[58]
  PIN dma_hrdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.680 4.000 849.280 ;
    END
  END dma_hrdata[59]
  PIN dma_hrdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END dma_hrdata[5]
  PIN dma_hrdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.720 4.000 851.320 ;
    END
  END dma_hrdata[60]
  PIN dma_hrdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.080 4.000 852.680 ;
    END
  END dma_hrdata[61]
  PIN dma_hrdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.120 4.000 854.720 ;
    END
  END dma_hrdata[62]
  PIN dma_hrdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 855.480 4.000 856.080 ;
    END
  END dma_hrdata[63]
  PIN dma_hrdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.160 4.000 754.760 ;
    END
  END dma_hrdata[6]
  PIN dma_hrdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 755.520 4.000 756.120 ;
    END
  END dma_hrdata[7]
  PIN dma_hrdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END dma_hrdata[8]
  PIN dma_hrdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 759.600 4.000 760.200 ;
    END
  END dma_hrdata[9]
  PIN dma_hreadyin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END dma_hreadyin
  PIN dma_hreadyout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 857.520 4.000 858.120 ;
    END
  END dma_hreadyout
  PIN dma_hresp
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 859.560 4.000 860.160 ;
    END
  END dma_hresp
  PIN dma_hsel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END dma_hsel
  PIN dma_hsize[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.800 4.000 617.400 ;
    END
  END dma_hsize[0]
  PIN dma_hsize[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.160 4.000 618.760 ;
    END
  END dma_hsize[1]
  PIN dma_hsize[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END dma_hsize[2]
  PIN dma_htrans[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END dma_htrans[0]
  PIN dma_htrans[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END dma_htrans[1]
  PIN dma_hwdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END dma_hwdata[0]
  PIN dma_hwdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 645.360 4.000 645.960 ;
    END
  END dma_hwdata[10]
  PIN dma_hwdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END dma_hwdata[11]
  PIN dma_hwdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END dma_hwdata[12]
  PIN dma_hwdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END dma_hwdata[13]
  PIN dma_hwdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END dma_hwdata[14]
  PIN dma_hwdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END dma_hwdata[15]
  PIN dma_hwdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END dma_hwdata[16]
  PIN dma_hwdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 657.600 4.000 658.200 ;
    END
  END dma_hwdata[17]
  PIN dma_hwdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END dma_hwdata[18]
  PIN dma_hwdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END dma_hwdata[19]
  PIN dma_hwdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END dma_hwdata[1]
  PIN dma_hwdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END dma_hwdata[20]
  PIN dma_hwdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 664.400 4.000 665.000 ;
    END
  END dma_hwdata[21]
  PIN dma_hwdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END dma_hwdata[22]
  PIN dma_hwdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END dma_hwdata[23]
  PIN dma_hwdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END dma_hwdata[24]
  PIN dma_hwdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END dma_hwdata[25]
  PIN dma_hwdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.920 4.000 674.520 ;
    END
  END dma_hwdata[26]
  PIN dma_hwdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.280 4.000 675.880 ;
    END
  END dma_hwdata[27]
  PIN dma_hwdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END dma_hwdata[28]
  PIN dma_hwdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END dma_hwdata[29]
  PIN dma_hwdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END dma_hwdata[2]
  PIN dma_hwdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END dma_hwdata[30]
  PIN dma_hwdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END dma_hwdata[31]
  PIN dma_hwdata[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END dma_hwdata[32]
  PIN dma_hwdata[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.160 4.000 686.760 ;
    END
  END dma_hwdata[33]
  PIN dma_hwdata[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END dma_hwdata[34]
  PIN dma_hwdata[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END dma_hwdata[35]
  PIN dma_hwdata[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END dma_hwdata[36]
  PIN dma_hwdata[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.960 4.000 693.560 ;
    END
  END dma_hwdata[37]
  PIN dma_hwdata[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END dma_hwdata[38]
  PIN dma_hwdata[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END dma_hwdata[39]
  PIN dma_hwdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END dma_hwdata[3]
  PIN dma_hwdata[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 698.400 4.000 699.000 ;
    END
  END dma_hwdata[40]
  PIN dma_hwdata[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END dma_hwdata[41]
  PIN dma_hwdata[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 702.480 4.000 703.080 ;
    END
  END dma_hwdata[42]
  PIN dma_hwdata[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END dma_hwdata[43]
  PIN dma_hwdata[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END dma_hwdata[44]
  PIN dma_hwdata[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END dma_hwdata[45]
  PIN dma_hwdata[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.280 4.000 709.880 ;
    END
  END dma_hwdata[46]
  PIN dma_hwdata[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END dma_hwdata[47]
  PIN dma_hwdata[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END dma_hwdata[48]
  PIN dma_hwdata[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.720 4.000 715.320 ;
    END
  END dma_hwdata[49]
  PIN dma_hwdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 634.480 4.000 635.080 ;
    END
  END dma_hwdata[4]
  PIN dma_hwdata[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END dma_hwdata[50]
  PIN dma_hwdata[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END dma_hwdata[51]
  PIN dma_hwdata[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.160 4.000 720.760 ;
    END
  END dma_hwdata[52]
  PIN dma_hwdata[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 721.520 4.000 722.120 ;
    END
  END dma_hwdata[53]
  PIN dma_hwdata[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 723.560 4.000 724.160 ;
    END
  END dma_hwdata[54]
  PIN dma_hwdata[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 725.600 4.000 726.200 ;
    END
  END dma_hwdata[55]
  PIN dma_hwdata[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.960 4.000 727.560 ;
    END
  END dma_hwdata[56]
  PIN dma_hwdata[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.000 4.000 729.600 ;
    END
  END dma_hwdata[57]
  PIN dma_hwdata[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END dma_hwdata[58]
  PIN dma_hwdata[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 732.400 4.000 733.000 ;
    END
  END dma_hwdata[59]
  PIN dma_hwdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END dma_hwdata[5]
  PIN dma_hwdata[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END dma_hwdata[60]
  PIN dma_hwdata[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END dma_hwdata[61]
  PIN dma_hwdata[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END dma_hwdata[62]
  PIN dma_hwdata[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.880 4.000 740.480 ;
    END
  END dma_hwdata[63]
  PIN dma_hwdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END dma_hwdata[6]
  PIN dma_hwdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END dma_hwdata[7]
  PIN dma_hwdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.280 4.000 641.880 ;
    END
  END dma_hwdata[8]
  PIN dma_hwdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END dma_hwdata[9]
  PIN dma_hwrite
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END dma_hwrite
  PIN extintsrc_req[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END extintsrc_req[0]
  PIN extintsrc_req[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END extintsrc_req[10]
  PIN extintsrc_req[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END extintsrc_req[11]
  PIN extintsrc_req[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END extintsrc_req[12]
  PIN extintsrc_req[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END extintsrc_req[13]
  PIN extintsrc_req[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END extintsrc_req[14]
  PIN extintsrc_req[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END extintsrc_req[15]
  PIN extintsrc_req[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END extintsrc_req[16]
  PIN extintsrc_req[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END extintsrc_req[17]
  PIN extintsrc_req[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END extintsrc_req[18]
  PIN extintsrc_req[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END extintsrc_req[19]
  PIN extintsrc_req[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END extintsrc_req[1]
  PIN extintsrc_req[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END extintsrc_req[20]
  PIN extintsrc_req[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END extintsrc_req[21]
  PIN extintsrc_req[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END extintsrc_req[22]
  PIN extintsrc_req[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END extintsrc_req[23]
  PIN extintsrc_req[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END extintsrc_req[24]
  PIN extintsrc_req[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END extintsrc_req[25]
  PIN extintsrc_req[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END extintsrc_req[26]
  PIN extintsrc_req[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END extintsrc_req[27]
  PIN extintsrc_req[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END extintsrc_req[28]
  PIN extintsrc_req[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END extintsrc_req[29]
  PIN extintsrc_req[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END extintsrc_req[2]
  PIN extintsrc_req[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END extintsrc_req[30]
  PIN extintsrc_req[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END extintsrc_req[3]
  PIN extintsrc_req[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END extintsrc_req[4]
  PIN extintsrc_req[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END extintsrc_req[5]
  PIN extintsrc_req[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END extintsrc_req[6]
  PIN extintsrc_req[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END extintsrc_req[7]
  PIN extintsrc_req[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END extintsrc_req[8]
  PIN extintsrc_req[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END extintsrc_req[9]
  PIN haddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END haddr[0]
  PIN haddr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END haddr[10]
  PIN haddr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END haddr[11]
  PIN haddr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END haddr[12]
  PIN haddr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END haddr[13]
  PIN haddr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END haddr[14]
  PIN haddr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END haddr[15]
  PIN haddr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END haddr[16]
  PIN haddr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END haddr[17]
  PIN haddr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END haddr[18]
  PIN haddr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END haddr[19]
  PIN haddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END haddr[1]
  PIN haddr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END haddr[20]
  PIN haddr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END haddr[21]
  PIN haddr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END haddr[22]
  PIN haddr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END haddr[23]
  PIN haddr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END haddr[24]
  PIN haddr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END haddr[25]
  PIN haddr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END haddr[26]
  PIN haddr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END haddr[27]
  PIN haddr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END haddr[28]
  PIN haddr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END haddr[29]
  PIN haddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END haddr[2]
  PIN haddr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END haddr[30]
  PIN haddr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END haddr[31]
  PIN haddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END haddr[3]
  PIN haddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END haddr[4]
  PIN haddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END haddr[5]
  PIN haddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END haddr[6]
  PIN haddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END haddr[7]
  PIN haddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END haddr[8]
  PIN haddr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END haddr[9]
  PIN hburst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END hburst[0]
  PIN hburst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END hburst[1]
  PIN hburst[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END hburst[2]
  PIN hmastlock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END hmastlock
  PIN hprot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END hprot[0]
  PIN hprot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END hprot[1]
  PIN hprot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END hprot[2]
  PIN hprot[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END hprot[3]
  PIN hrdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END hrdata[0]
  PIN hrdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END hrdata[10]
  PIN hrdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END hrdata[11]
  PIN hrdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END hrdata[12]
  PIN hrdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END hrdata[13]
  PIN hrdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END hrdata[14]
  PIN hrdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END hrdata[15]
  PIN hrdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END hrdata[16]
  PIN hrdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END hrdata[17]
  PIN hrdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END hrdata[18]
  PIN hrdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END hrdata[19]
  PIN hrdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END hrdata[1]
  PIN hrdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END hrdata[20]
  PIN hrdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END hrdata[21]
  PIN hrdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END hrdata[22]
  PIN hrdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END hrdata[23]
  PIN hrdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END hrdata[24]
  PIN hrdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END hrdata[25]
  PIN hrdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END hrdata[26]
  PIN hrdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 0.000 510.510 4.000 ;
    END
  END hrdata[27]
  PIN hrdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END hrdata[28]
  PIN hrdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END hrdata[29]
  PIN hrdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END hrdata[2]
  PIN hrdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END hrdata[30]
  PIN hrdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END hrdata[31]
  PIN hrdata[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END hrdata[32]
  PIN hrdata[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END hrdata[33]
  PIN hrdata[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END hrdata[34]
  PIN hrdata[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END hrdata[35]
  PIN hrdata[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END hrdata[36]
  PIN hrdata[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END hrdata[37]
  PIN hrdata[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END hrdata[38]
  PIN hrdata[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END hrdata[39]
  PIN hrdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END hrdata[3]
  PIN hrdata[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END hrdata[40]
  PIN hrdata[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END hrdata[41]
  PIN hrdata[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END hrdata[42]
  PIN hrdata[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END hrdata[43]
  PIN hrdata[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END hrdata[44]
  PIN hrdata[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END hrdata[45]
  PIN hrdata[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END hrdata[46]
  PIN hrdata[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END hrdata[47]
  PIN hrdata[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END hrdata[48]
  PIN hrdata[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END hrdata[49]
  PIN hrdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END hrdata[4]
  PIN hrdata[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END hrdata[50]
  PIN hrdata[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END hrdata[51]
  PIN hrdata[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 0.000 645.750 4.000 ;
    END
  END hrdata[52]
  PIN hrdata[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END hrdata[53]
  PIN hrdata[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END hrdata[54]
  PIN hrdata[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END hrdata[55]
  PIN hrdata[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END hrdata[56]
  PIN hrdata[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 0.000 672.430 4.000 ;
    END
  END hrdata[57]
  PIN hrdata[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 0.000 677.950 4.000 ;
    END
  END hrdata[58]
  PIN hrdata[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END hrdata[59]
  PIN hrdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END hrdata[5]
  PIN hrdata[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END hrdata[60]
  PIN hrdata[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 0.000 694.050 4.000 ;
    END
  END hrdata[61]
  PIN hrdata[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END hrdata[62]
  PIN hrdata[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 0.000 705.090 4.000 ;
    END
  END hrdata[63]
  PIN hrdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END hrdata[6]
  PIN hrdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END hrdata[7]
  PIN hrdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END hrdata[8]
  PIN hrdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END hrdata[9]
  PIN hready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END hready
  PIN hresp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END hresp
  PIN hsize[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END hsize[0]
  PIN hsize[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END hsize[1]
  PIN hsize[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END hsize[2]
  PIN htrans[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END htrans[0]
  PIN htrans[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END htrans[1]
  PIN hwrite
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END hwrite
  PIN i_cpu_halt_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1300.200 4.000 1300.800 ;
    END
  END i_cpu_halt_req
  PIN i_cpu_run_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1307.680 4.000 1308.280 ;
    END
  END i_cpu_run_req
  PIN ic_data_ext_in_pkt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1039.760 4.000 1040.360 ;
    END
  END ic_data_ext_in_pkt[0]
  PIN ic_data_ext_in_pkt[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END ic_data_ext_in_pkt[10]
  PIN ic_data_ext_in_pkt[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1059.480 4.000 1060.080 ;
    END
  END ic_data_ext_in_pkt[11]
  PIN ic_data_ext_in_pkt[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END ic_data_ext_in_pkt[12]
  PIN ic_data_ext_in_pkt[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1062.880 4.000 1063.480 ;
    END
  END ic_data_ext_in_pkt[13]
  PIN ic_data_ext_in_pkt[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.920 4.000 1065.520 ;
    END
  END ic_data_ext_in_pkt[14]
  PIN ic_data_ext_in_pkt[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.280 4.000 1066.880 ;
    END
  END ic_data_ext_in_pkt[15]
  PIN ic_data_ext_in_pkt[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1068.320 4.000 1068.920 ;
    END
  END ic_data_ext_in_pkt[16]
  PIN ic_data_ext_in_pkt[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1070.360 4.000 1070.960 ;
    END
  END ic_data_ext_in_pkt[17]
  PIN ic_data_ext_in_pkt[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.720 4.000 1072.320 ;
    END
  END ic_data_ext_in_pkt[18]
  PIN ic_data_ext_in_pkt[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1073.760 4.000 1074.360 ;
    END
  END ic_data_ext_in_pkt[19]
  PIN ic_data_ext_in_pkt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.800 4.000 1042.400 ;
    END
  END ic_data_ext_in_pkt[1]
  PIN ic_data_ext_in_pkt[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.120 4.000 1075.720 ;
    END
  END ic_data_ext_in_pkt[20]
  PIN ic_data_ext_in_pkt[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.160 4.000 1077.760 ;
    END
  END ic_data_ext_in_pkt[21]
  PIN ic_data_ext_in_pkt[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1079.200 4.000 1079.800 ;
    END
  END ic_data_ext_in_pkt[22]
  PIN ic_data_ext_in_pkt[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1080.560 4.000 1081.160 ;
    END
  END ic_data_ext_in_pkt[23]
  PIN ic_data_ext_in_pkt[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1082.600 4.000 1083.200 ;
    END
  END ic_data_ext_in_pkt[24]
  PIN ic_data_ext_in_pkt[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END ic_data_ext_in_pkt[25]
  PIN ic_data_ext_in_pkt[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1086.000 4.000 1086.600 ;
    END
  END ic_data_ext_in_pkt[26]
  PIN ic_data_ext_in_pkt[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END ic_data_ext_in_pkt[27]
  PIN ic_data_ext_in_pkt[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1089.400 4.000 1090.000 ;
    END
  END ic_data_ext_in_pkt[28]
  PIN ic_data_ext_in_pkt[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END ic_data_ext_in_pkt[29]
  PIN ic_data_ext_in_pkt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.160 4.000 1043.760 ;
    END
  END ic_data_ext_in_pkt[2]
  PIN ic_data_ext_in_pkt[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1093.480 4.000 1094.080 ;
    END
  END ic_data_ext_in_pkt[30]
  PIN ic_data_ext_in_pkt[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END ic_data_ext_in_pkt[31]
  PIN ic_data_ext_in_pkt[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.880 4.000 1097.480 ;
    END
  END ic_data_ext_in_pkt[32]
  PIN ic_data_ext_in_pkt[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.920 4.000 1099.520 ;
    END
  END ic_data_ext_in_pkt[33]
  PIN ic_data_ext_in_pkt[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1100.280 4.000 1100.880 ;
    END
  END ic_data_ext_in_pkt[34]
  PIN ic_data_ext_in_pkt[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1102.320 4.000 1102.920 ;
    END
  END ic_data_ext_in_pkt[35]
  PIN ic_data_ext_in_pkt[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1103.680 4.000 1104.280 ;
    END
  END ic_data_ext_in_pkt[36]
  PIN ic_data_ext_in_pkt[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.720 4.000 1106.320 ;
    END
  END ic_data_ext_in_pkt[37]
  PIN ic_data_ext_in_pkt[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1107.760 4.000 1108.360 ;
    END
  END ic_data_ext_in_pkt[38]
  PIN ic_data_ext_in_pkt[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.120 4.000 1109.720 ;
    END
  END ic_data_ext_in_pkt[39]
  PIN ic_data_ext_in_pkt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.200 4.000 1045.800 ;
    END
  END ic_data_ext_in_pkt[3]
  PIN ic_data_ext_in_pkt[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.160 4.000 1111.760 ;
    END
  END ic_data_ext_in_pkt[40]
  PIN ic_data_ext_in_pkt[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1113.200 4.000 1113.800 ;
    END
  END ic_data_ext_in_pkt[41]
  PIN ic_data_ext_in_pkt[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1114.560 4.000 1115.160 ;
    END
  END ic_data_ext_in_pkt[42]
  PIN ic_data_ext_in_pkt[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1116.600 4.000 1117.200 ;
    END
  END ic_data_ext_in_pkt[43]
  PIN ic_data_ext_in_pkt[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1117.960 4.000 1118.560 ;
    END
  END ic_data_ext_in_pkt[44]
  PIN ic_data_ext_in_pkt[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.000 4.000 1120.600 ;
    END
  END ic_data_ext_in_pkt[45]
  PIN ic_data_ext_in_pkt[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END ic_data_ext_in_pkt[46]
  PIN ic_data_ext_in_pkt[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1123.400 4.000 1124.000 ;
    END
  END ic_data_ext_in_pkt[47]
  PIN ic_data_ext_in_pkt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1046.560 4.000 1047.160 ;
    END
  END ic_data_ext_in_pkt[4]
  PIN ic_data_ext_in_pkt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1048.600 4.000 1049.200 ;
    END
  END ic_data_ext_in_pkt[5]
  PIN ic_data_ext_in_pkt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END ic_data_ext_in_pkt[6]
  PIN ic_data_ext_in_pkt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1052.000 4.000 1052.600 ;
    END
  END ic_data_ext_in_pkt[7]
  PIN ic_data_ext_in_pkt[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END ic_data_ext_in_pkt[8]
  PIN ic_data_ext_in_pkt[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.080 4.000 1056.680 ;
    END
  END ic_data_ext_in_pkt[9]
  PIN ic_tag_ext_in_pkt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1125.440 4.000 1126.040 ;
    END
  END ic_tag_ext_in_pkt[0]
  PIN ic_tag_ext_in_pkt[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1143.120 4.000 1143.720 ;
    END
  END ic_tag_ext_in_pkt[10]
  PIN ic_tag_ext_in_pkt[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.160 4.000 1145.760 ;
    END
  END ic_tag_ext_in_pkt[11]
  PIN ic_tag_ext_in_pkt[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1147.200 4.000 1147.800 ;
    END
  END ic_tag_ext_in_pkt[12]
  PIN ic_tag_ext_in_pkt[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1148.560 4.000 1149.160 ;
    END
  END ic_tag_ext_in_pkt[13]
  PIN ic_tag_ext_in_pkt[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1150.600 4.000 1151.200 ;
    END
  END ic_tag_ext_in_pkt[14]
  PIN ic_tag_ext_in_pkt[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1151.960 4.000 1152.560 ;
    END
  END ic_tag_ext_in_pkt[15]
  PIN ic_tag_ext_in_pkt[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1154.000 4.000 1154.600 ;
    END
  END ic_tag_ext_in_pkt[16]
  PIN ic_tag_ext_in_pkt[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END ic_tag_ext_in_pkt[17]
  PIN ic_tag_ext_in_pkt[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1157.400 4.000 1158.000 ;
    END
  END ic_tag_ext_in_pkt[18]
  PIN ic_tag_ext_in_pkt[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1159.440 4.000 1160.040 ;
    END
  END ic_tag_ext_in_pkt[19]
  PIN ic_tag_ext_in_pkt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1127.480 4.000 1128.080 ;
    END
  END ic_tag_ext_in_pkt[1]
  PIN ic_tag_ext_in_pkt[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1161.480 4.000 1162.080 ;
    END
  END ic_tag_ext_in_pkt[20]
  PIN ic_tag_ext_in_pkt[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END ic_tag_ext_in_pkt[21]
  PIN ic_tag_ext_in_pkt[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1164.880 4.000 1165.480 ;
    END
  END ic_tag_ext_in_pkt[22]
  PIN ic_tag_ext_in_pkt[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END ic_tag_ext_in_pkt[23]
  PIN ic_tag_ext_in_pkt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END ic_tag_ext_in_pkt[2]
  PIN ic_tag_ext_in_pkt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1130.880 4.000 1131.480 ;
    END
  END ic_tag_ext_in_pkt[3]
  PIN ic_tag_ext_in_pkt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.920 4.000 1133.520 ;
    END
  END ic_tag_ext_in_pkt[4]
  PIN ic_tag_ext_in_pkt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1134.280 4.000 1134.880 ;
    END
  END ic_tag_ext_in_pkt[5]
  PIN ic_tag_ext_in_pkt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1136.320 4.000 1136.920 ;
    END
  END ic_tag_ext_in_pkt[6]
  PIN ic_tag_ext_in_pkt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1137.680 4.000 1138.280 ;
    END
  END ic_tag_ext_in_pkt[7]
  PIN ic_tag_ext_in_pkt[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.720 4.000 1140.320 ;
    END
  END ic_tag_ext_in_pkt[8]
  PIN ic_tag_ext_in_pkt[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.760 4.000 1142.360 ;
    END
  END ic_tag_ext_in_pkt[9]
  PIN iccm_ext_in_pkt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 954.080 4.000 954.680 ;
    END
  END iccm_ext_in_pkt[0]
  PIN iccm_ext_in_pkt[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.760 4.000 972.360 ;
    END
  END iccm_ext_in_pkt[10]
  PIN iccm_ext_in_pkt[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 973.800 4.000 974.400 ;
    END
  END iccm_ext_in_pkt[11]
  PIN iccm_ext_in_pkt[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.160 4.000 975.760 ;
    END
  END iccm_ext_in_pkt[12]
  PIN iccm_ext_in_pkt[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.200 4.000 977.800 ;
    END
  END iccm_ext_in_pkt[13]
  PIN iccm_ext_in_pkt[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END iccm_ext_in_pkt[14]
  PIN iccm_ext_in_pkt[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END iccm_ext_in_pkt[15]
  PIN iccm_ext_in_pkt[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 982.640 4.000 983.240 ;
    END
  END iccm_ext_in_pkt[16]
  PIN iccm_ext_in_pkt[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 984.680 4.000 985.280 ;
    END
  END iccm_ext_in_pkt[17]
  PIN iccm_ext_in_pkt[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END iccm_ext_in_pkt[18]
  PIN iccm_ext_in_pkt[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 988.080 4.000 988.680 ;
    END
  END iccm_ext_in_pkt[19]
  PIN iccm_ext_in_pkt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 956.120 4.000 956.720 ;
    END
  END iccm_ext_in_pkt[1]
  PIN iccm_ext_in_pkt[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END iccm_ext_in_pkt[20]
  PIN iccm_ext_in_pkt[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 991.480 4.000 992.080 ;
    END
  END iccm_ext_in_pkt[21]
  PIN iccm_ext_in_pkt[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 993.520 4.000 994.120 ;
    END
  END iccm_ext_in_pkt[22]
  PIN iccm_ext_in_pkt[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.880 4.000 995.480 ;
    END
  END iccm_ext_in_pkt[23]
  PIN iccm_ext_in_pkt[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.920 4.000 997.520 ;
    END
  END iccm_ext_in_pkt[24]
  PIN iccm_ext_in_pkt[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 998.960 4.000 999.560 ;
    END
  END iccm_ext_in_pkt[25]
  PIN iccm_ext_in_pkt[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1000.320 4.000 1000.920 ;
    END
  END iccm_ext_in_pkt[26]
  PIN iccm_ext_in_pkt[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1002.360 4.000 1002.960 ;
    END
  END iccm_ext_in_pkt[27]
  PIN iccm_ext_in_pkt[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.720 4.000 1004.320 ;
    END
  END iccm_ext_in_pkt[28]
  PIN iccm_ext_in_pkt[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1005.760 4.000 1006.360 ;
    END
  END iccm_ext_in_pkt[29]
  PIN iccm_ext_in_pkt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 957.480 4.000 958.080 ;
    END
  END iccm_ext_in_pkt[2]
  PIN iccm_ext_in_pkt[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.800 4.000 1008.400 ;
    END
  END iccm_ext_in_pkt[30]
  PIN iccm_ext_in_pkt[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.160 4.000 1009.760 ;
    END
  END iccm_ext_in_pkt[31]
  PIN iccm_ext_in_pkt[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.200 4.000 1011.800 ;
    END
  END iccm_ext_in_pkt[32]
  PIN iccm_ext_in_pkt[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END iccm_ext_in_pkt[33]
  PIN iccm_ext_in_pkt[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1014.600 4.000 1015.200 ;
    END
  END iccm_ext_in_pkt[34]
  PIN iccm_ext_in_pkt[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1016.640 4.000 1017.240 ;
    END
  END iccm_ext_in_pkt[35]
  PIN iccm_ext_in_pkt[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.000 4.000 1018.600 ;
    END
  END iccm_ext_in_pkt[36]
  PIN iccm_ext_in_pkt[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END iccm_ext_in_pkt[37]
  PIN iccm_ext_in_pkt[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1022.080 4.000 1022.680 ;
    END
  END iccm_ext_in_pkt[38]
  PIN iccm_ext_in_pkt[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1023.440 4.000 1024.040 ;
    END
  END iccm_ext_in_pkt[39]
  PIN iccm_ext_in_pkt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 959.520 4.000 960.120 ;
    END
  END iccm_ext_in_pkt[3]
  PIN iccm_ext_in_pkt[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1025.480 4.000 1026.080 ;
    END
  END iccm_ext_in_pkt[40]
  PIN iccm_ext_in_pkt[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1027.520 4.000 1028.120 ;
    END
  END iccm_ext_in_pkt[41]
  PIN iccm_ext_in_pkt[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1028.880 4.000 1029.480 ;
    END
  END iccm_ext_in_pkt[42]
  PIN iccm_ext_in_pkt[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.920 4.000 1031.520 ;
    END
  END iccm_ext_in_pkt[43]
  PIN iccm_ext_in_pkt[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.280 4.000 1032.880 ;
    END
  END iccm_ext_in_pkt[44]
  PIN iccm_ext_in_pkt[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1034.320 4.000 1034.920 ;
    END
  END iccm_ext_in_pkt[45]
  PIN iccm_ext_in_pkt[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END iccm_ext_in_pkt[46]
  PIN iccm_ext_in_pkt[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.720 4.000 1038.320 ;
    END
  END iccm_ext_in_pkt[47]
  PIN iccm_ext_in_pkt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.880 4.000 961.480 ;
    END
  END iccm_ext_in_pkt[4]
  PIN iccm_ext_in_pkt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.920 4.000 963.520 ;
    END
  END iccm_ext_in_pkt[5]
  PIN iccm_ext_in_pkt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.960 4.000 965.560 ;
    END
  END iccm_ext_in_pkt[6]
  PIN iccm_ext_in_pkt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 966.320 4.000 966.920 ;
    END
  END iccm_ext_in_pkt[7]
  PIN iccm_ext_in_pkt[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 968.360 4.000 968.960 ;
    END
  END iccm_ext_in_pkt[8]
  PIN iccm_ext_in_pkt[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 970.400 4.000 971.000 ;
    END
  END iccm_ext_in_pkt[9]
  PIN ifu_bus_clk_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.960 4.000 863.560 ;
    END
  END ifu_bus_clk_en
  PIN jtag_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1184.600 4.000 1185.200 ;
    END
  END jtag_id[0]
  PIN jtag_id[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1202.280 4.000 1202.880 ;
    END
  END jtag_id[10]
  PIN jtag_id[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1204.320 4.000 1204.920 ;
    END
  END jtag_id[11]
  PIN jtag_id[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1205.680 4.000 1206.280 ;
    END
  END jtag_id[12]
  PIN jtag_id[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.720 4.000 1208.320 ;
    END
  END jtag_id[13]
  PIN jtag_id[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1209.080 4.000 1209.680 ;
    END
  END jtag_id[14]
  PIN jtag_id[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1211.120 4.000 1211.720 ;
    END
  END jtag_id[15]
  PIN jtag_id[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.160 4.000 1213.760 ;
    END
  END jtag_id[16]
  PIN jtag_id[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1214.520 4.000 1215.120 ;
    END
  END jtag_id[17]
  PIN jtag_id[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1216.560 4.000 1217.160 ;
    END
  END jtag_id[18]
  PIN jtag_id[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1218.600 4.000 1219.200 ;
    END
  END jtag_id[19]
  PIN jtag_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1185.960 4.000 1186.560 ;
    END
  END jtag_id[1]
  PIN jtag_id[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1219.960 4.000 1220.560 ;
    END
  END jtag_id[20]
  PIN jtag_id[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1222.000 4.000 1222.600 ;
    END
  END jtag_id[21]
  PIN jtag_id[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1223.360 4.000 1223.960 ;
    END
  END jtag_id[22]
  PIN jtag_id[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1225.400 4.000 1226.000 ;
    END
  END jtag_id[23]
  PIN jtag_id[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END jtag_id[24]
  PIN jtag_id[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1228.800 4.000 1229.400 ;
    END
  END jtag_id[25]
  PIN jtag_id[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.840 4.000 1231.440 ;
    END
  END jtag_id[26]
  PIN jtag_id[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1232.880 4.000 1233.480 ;
    END
  END jtag_id[27]
  PIN jtag_id[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1234.240 4.000 1234.840 ;
    END
  END jtag_id[28]
  PIN jtag_id[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.280 4.000 1236.880 ;
    END
  END jtag_id[29]
  PIN jtag_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1188.000 4.000 1188.600 ;
    END
  END jtag_id[2]
  PIN jtag_id[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1237.640 4.000 1238.240 ;
    END
  END jtag_id[30]
  PIN jtag_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.040 4.000 1190.640 ;
    END
  END jtag_id[3]
  PIN jtag_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1191.400 4.000 1192.000 ;
    END
  END jtag_id[4]
  PIN jtag_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END jtag_id[5]
  PIN jtag_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.800 4.000 1195.400 ;
    END
  END jtag_id[6]
  PIN jtag_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1196.840 4.000 1197.440 ;
    END
  END jtag_id[7]
  PIN jtag_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1198.880 4.000 1199.480 ;
    END
  END jtag_id[8]
  PIN jtag_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.240 4.000 1200.840 ;
    END
  END jtag_id[9]
  PIN jtag_tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1175.760 4.000 1176.360 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.160 4.000 1179.760 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1182.560 4.000 1183.160 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1177.120 4.000 1177.720 ;
    END
  END jtag_tms
  PIN jtag_trst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1180.520 4.000 1181.120 ;
    END
  END jtag_trst_n
  PIN lsu_bus_clk_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.920 4.000 861.520 ;
    END
  END lsu_bus_clk_en
  PIN lsu_haddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END lsu_haddr[0]
  PIN lsu_haddr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END lsu_haddr[10]
  PIN lsu_haddr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END lsu_haddr[11]
  PIN lsu_haddr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END lsu_haddr[12]
  PIN lsu_haddr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END lsu_haddr[13]
  PIN lsu_haddr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END lsu_haddr[14]
  PIN lsu_haddr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END lsu_haddr[15]
  PIN lsu_haddr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END lsu_haddr[16]
  PIN lsu_haddr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END lsu_haddr[17]
  PIN lsu_haddr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END lsu_haddr[18]
  PIN lsu_haddr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END lsu_haddr[19]
  PIN lsu_haddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END lsu_haddr[1]
  PIN lsu_haddr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END lsu_haddr[20]
  PIN lsu_haddr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END lsu_haddr[21]
  PIN lsu_haddr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END lsu_haddr[22]
  PIN lsu_haddr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END lsu_haddr[23]
  PIN lsu_haddr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END lsu_haddr[24]
  PIN lsu_haddr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 4.000 ;
    END
  END lsu_haddr[25]
  PIN lsu_haddr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END lsu_haddr[26]
  PIN lsu_haddr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END lsu_haddr[27]
  PIN lsu_haddr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END lsu_haddr[28]
  PIN lsu_haddr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END lsu_haddr[29]
  PIN lsu_haddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END lsu_haddr[2]
  PIN lsu_haddr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END lsu_haddr[30]
  PIN lsu_haddr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END lsu_haddr[31]
  PIN lsu_haddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END lsu_haddr[3]
  PIN lsu_haddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END lsu_haddr[4]
  PIN lsu_haddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END lsu_haddr[5]
  PIN lsu_haddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END lsu_haddr[6]
  PIN lsu_haddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END lsu_haddr[7]
  PIN lsu_haddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END lsu_haddr[8]
  PIN lsu_haddr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END lsu_haddr[9]
  PIN lsu_hburst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END lsu_hburst[0]
  PIN lsu_hburst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END lsu_hburst[1]
  PIN lsu_hburst[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END lsu_hburst[2]
  PIN lsu_hmastlock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END lsu_hmastlock
  PIN lsu_hprot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END lsu_hprot[0]
  PIN lsu_hprot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END lsu_hprot[1]
  PIN lsu_hprot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END lsu_hprot[2]
  PIN lsu_hprot[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END lsu_hprot[3]
  PIN lsu_hrdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END lsu_hrdata[0]
  PIN lsu_hrdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 0.000 764.430 4.000 ;
    END
  END lsu_hrdata[10]
  PIN lsu_hrdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END lsu_hrdata[11]
  PIN lsu_hrdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 0.000 775.470 4.000 ;
    END
  END lsu_hrdata[12]
  PIN lsu_hrdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END lsu_hrdata[13]
  PIN lsu_hrdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END lsu_hrdata[14]
  PIN lsu_hrdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 0.000 791.570 4.000 ;
    END
  END lsu_hrdata[15]
  PIN lsu_hrdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 4.000 ;
    END
  END lsu_hrdata[16]
  PIN lsu_hrdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END lsu_hrdata[17]
  PIN lsu_hrdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 0.000 807.670 4.000 ;
    END
  END lsu_hrdata[18]
  PIN lsu_hrdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.910 0.000 813.190 4.000 ;
    END
  END lsu_hrdata[19]
  PIN lsu_hrdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END lsu_hrdata[1]
  PIN lsu_hrdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 4.000 ;
    END
  END lsu_hrdata[20]
  PIN lsu_hrdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.490 0.000 823.770 4.000 ;
    END
  END lsu_hrdata[21]
  PIN lsu_hrdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 0.000 829.290 4.000 ;
    END
  END lsu_hrdata[22]
  PIN lsu_hrdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 0.000 834.810 4.000 ;
    END
  END lsu_hrdata[23]
  PIN lsu_hrdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 0.000 840.330 4.000 ;
    END
  END lsu_hrdata[24]
  PIN lsu_hrdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 0.000 845.390 4.000 ;
    END
  END lsu_hrdata[25]
  PIN lsu_hrdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 0.000 850.910 4.000 ;
    END
  END lsu_hrdata[26]
  PIN lsu_hrdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 0.000 856.430 4.000 ;
    END
  END lsu_hrdata[27]
  PIN lsu_hrdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 0.000 861.950 4.000 ;
    END
  END lsu_hrdata[28]
  PIN lsu_hrdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 0.000 867.010 4.000 ;
    END
  END lsu_hrdata[29]
  PIN lsu_hrdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END lsu_hrdata[2]
  PIN lsu_hrdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END lsu_hrdata[30]
  PIN lsu_hrdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 0.000 878.050 4.000 ;
    END
  END lsu_hrdata[31]
  PIN lsu_hrdata[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 0.000 883.570 4.000 ;
    END
  END lsu_hrdata[32]
  PIN lsu_hrdata[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END lsu_hrdata[33]
  PIN lsu_hrdata[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 0.000 894.150 4.000 ;
    END
  END lsu_hrdata[34]
  PIN lsu_hrdata[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END lsu_hrdata[35]
  PIN lsu_hrdata[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END lsu_hrdata[36]
  PIN lsu_hrdata[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.970 0.000 910.250 4.000 ;
    END
  END lsu_hrdata[37]
  PIN lsu_hrdata[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.490 0.000 915.770 4.000 ;
    END
  END lsu_hrdata[38]
  PIN lsu_hrdata[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END lsu_hrdata[39]
  PIN lsu_hrdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 0.000 726.710 4.000 ;
    END
  END lsu_hrdata[3]
  PIN lsu_hrdata[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.530 0.000 926.810 4.000 ;
    END
  END lsu_hrdata[40]
  PIN lsu_hrdata[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 0.000 931.870 4.000 ;
    END
  END lsu_hrdata[41]
  PIN lsu_hrdata[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END lsu_hrdata[42]
  PIN lsu_hrdata[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 0.000 942.910 4.000 ;
    END
  END lsu_hrdata[43]
  PIN lsu_hrdata[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 0.000 948.430 4.000 ;
    END
  END lsu_hrdata[44]
  PIN lsu_hrdata[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END lsu_hrdata[45]
  PIN lsu_hrdata[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 0.000 959.010 4.000 ;
    END
  END lsu_hrdata[46]
  PIN lsu_hrdata[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.250 0.000 964.530 4.000 ;
    END
  END lsu_hrdata[47]
  PIN lsu_hrdata[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 0.000 970.050 4.000 ;
    END
  END lsu_hrdata[48]
  PIN lsu_hrdata[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.830 0.000 975.110 4.000 ;
    END
  END lsu_hrdata[49]
  PIN lsu_hrdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 0.000 732.230 4.000 ;
    END
  END lsu_hrdata[4]
  PIN lsu_hrdata[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 0.000 980.630 4.000 ;
    END
  END lsu_hrdata[50]
  PIN lsu_hrdata[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.870 0.000 986.150 4.000 ;
    END
  END lsu_hrdata[51]
  PIN lsu_hrdata[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 0.000 991.670 4.000 ;
    END
  END lsu_hrdata[52]
  PIN lsu_hrdata[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 0.000 996.730 4.000 ;
    END
  END lsu_hrdata[53]
  PIN lsu_hrdata[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.970 0.000 1002.250 4.000 ;
    END
  END lsu_hrdata[54]
  PIN lsu_hrdata[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.490 0.000 1007.770 4.000 ;
    END
  END lsu_hrdata[55]
  PIN lsu_hrdata[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 0.000 1013.290 4.000 ;
    END
  END lsu_hrdata[56]
  PIN lsu_hrdata[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.070 0.000 1018.350 4.000 ;
    END
  END lsu_hrdata[57]
  PIN lsu_hrdata[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.590 0.000 1023.870 4.000 ;
    END
  END lsu_hrdata[58]
  PIN lsu_hrdata[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 0.000 1029.390 4.000 ;
    END
  END lsu_hrdata[59]
  PIN lsu_hrdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END lsu_hrdata[5]
  PIN lsu_hrdata[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.630 0.000 1034.910 4.000 ;
    END
  END lsu_hrdata[60]
  PIN lsu_hrdata[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.690 0.000 1039.970 4.000 ;
    END
  END lsu_hrdata[61]
  PIN lsu_hrdata[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.210 0.000 1045.490 4.000 ;
    END
  END lsu_hrdata[62]
  PIN lsu_hrdata[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.730 0.000 1051.010 4.000 ;
    END
  END lsu_hrdata[63]
  PIN lsu_hrdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 0.000 742.810 4.000 ;
    END
  END lsu_hrdata[6]
  PIN lsu_hrdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END lsu_hrdata[7]
  PIN lsu_hrdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END lsu_hrdata[8]
  PIN lsu_hrdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.630 0.000 758.910 4.000 ;
    END
  END lsu_hrdata[9]
  PIN lsu_hready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END lsu_hready
  PIN lsu_hresp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END lsu_hresp
  PIN lsu_hsize[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END lsu_hsize[0]
  PIN lsu_hsize[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END lsu_hsize[1]
  PIN lsu_hsize[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END lsu_hsize[2]
  PIN lsu_htrans[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END lsu_htrans[0]
  PIN lsu_htrans[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END lsu_htrans[1]
  PIN lsu_hwdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END lsu_hwdata[0]
  PIN lsu_hwdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 0.000 1110.350 4.000 ;
    END
  END lsu_hwdata[10]
  PIN lsu_hwdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.590 0.000 1115.870 4.000 ;
    END
  END lsu_hwdata[11]
  PIN lsu_hwdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 0.000 1121.390 4.000 ;
    END
  END lsu_hwdata[12]
  PIN lsu_hwdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.170 0.000 1126.450 4.000 ;
    END
  END lsu_hwdata[13]
  PIN lsu_hwdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.690 0.000 1131.970 4.000 ;
    END
  END lsu_hwdata[14]
  PIN lsu_hwdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 0.000 1137.490 4.000 ;
    END
  END lsu_hwdata[15]
  PIN lsu_hwdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.730 0.000 1143.010 4.000 ;
    END
  END lsu_hwdata[16]
  PIN lsu_hwdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.790 0.000 1148.070 4.000 ;
    END
  END lsu_hwdata[17]
  PIN lsu_hwdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.310 0.000 1153.590 4.000 ;
    END
  END lsu_hwdata[18]
  PIN lsu_hwdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.830 0.000 1159.110 4.000 ;
    END
  END lsu_hwdata[19]
  PIN lsu_hwdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.310 0.000 1061.590 4.000 ;
    END
  END lsu_hwdata[1]
  PIN lsu_hwdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END lsu_hwdata[20]
  PIN lsu_hwdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.410 0.000 1169.690 4.000 ;
    END
  END lsu_hwdata[21]
  PIN lsu_hwdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.930 0.000 1175.210 4.000 ;
    END
  END lsu_hwdata[22]
  PIN lsu_hwdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.450 0.000 1180.730 4.000 ;
    END
  END lsu_hwdata[23]
  PIN lsu_hwdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.970 0.000 1186.250 4.000 ;
    END
  END lsu_hwdata[24]
  PIN lsu_hwdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.030 0.000 1191.310 4.000 ;
    END
  END lsu_hwdata[25]
  PIN lsu_hwdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.550 0.000 1196.830 4.000 ;
    END
  END lsu_hwdata[26]
  PIN lsu_hwdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.070 0.000 1202.350 4.000 ;
    END
  END lsu_hwdata[27]
  PIN lsu_hwdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END lsu_hwdata[28]
  PIN lsu_hwdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.650 0.000 1212.930 4.000 ;
    END
  END lsu_hwdata[29]
  PIN lsu_hwdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.830 0.000 1067.110 4.000 ;
    END
  END lsu_hwdata[2]
  PIN lsu_hwdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 0.000 1218.450 4.000 ;
    END
  END lsu_hwdata[30]
  PIN lsu_hwdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 0.000 1223.970 4.000 ;
    END
  END lsu_hwdata[31]
  PIN lsu_hwdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.210 0.000 1229.490 4.000 ;
    END
  END lsu_hwdata[32]
  PIN lsu_hwdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.270 0.000 1234.550 4.000 ;
    END
  END lsu_hwdata[33]
  PIN lsu_hwdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 0.000 1240.070 4.000 ;
    END
  END lsu_hwdata[34]
  PIN lsu_hwdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.310 0.000 1245.590 4.000 ;
    END
  END lsu_hwdata[35]
  PIN lsu_hwdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.830 0.000 1251.110 4.000 ;
    END
  END lsu_hwdata[36]
  PIN lsu_hwdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 0.000 1256.170 4.000 ;
    END
  END lsu_hwdata[37]
  PIN lsu_hwdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.410 0.000 1261.690 4.000 ;
    END
  END lsu_hwdata[38]
  PIN lsu_hwdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.930 0.000 1267.210 4.000 ;
    END
  END lsu_hwdata[39]
  PIN lsu_hwdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END lsu_hwdata[3]
  PIN lsu_hwdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.450 0.000 1272.730 4.000 ;
    END
  END lsu_hwdata[40]
  PIN lsu_hwdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.510 0.000 1277.790 4.000 ;
    END
  END lsu_hwdata[41]
  PIN lsu_hwdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.030 0.000 1283.310 4.000 ;
    END
  END lsu_hwdata[42]
  PIN lsu_hwdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.550 0.000 1288.830 4.000 ;
    END
  END lsu_hwdata[43]
  PIN lsu_hwdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.070 0.000 1294.350 4.000 ;
    END
  END lsu_hwdata[44]
  PIN lsu_hwdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.130 0.000 1299.410 4.000 ;
    END
  END lsu_hwdata[45]
  PIN lsu_hwdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.650 0.000 1304.930 4.000 ;
    END
  END lsu_hwdata[46]
  PIN lsu_hwdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.170 0.000 1310.450 4.000 ;
    END
  END lsu_hwdata[47]
  PIN lsu_hwdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.690 0.000 1315.970 4.000 ;
    END
  END lsu_hwdata[48]
  PIN lsu_hwdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.750 0.000 1321.030 4.000 ;
    END
  END lsu_hwdata[49]
  PIN lsu_hwdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.870 0.000 1078.150 4.000 ;
    END
  END lsu_hwdata[4]
  PIN lsu_hwdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.270 0.000 1326.550 4.000 ;
    END
  END lsu_hwdata[50]
  PIN lsu_hwdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.790 0.000 1332.070 4.000 ;
    END
  END lsu_hwdata[51]
  PIN lsu_hwdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.310 0.000 1337.590 4.000 ;
    END
  END lsu_hwdata[52]
  PIN lsu_hwdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 0.000 1342.650 4.000 ;
    END
  END lsu_hwdata[53]
  PIN lsu_hwdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1347.890 0.000 1348.170 4.000 ;
    END
  END lsu_hwdata[54]
  PIN lsu_hwdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1353.410 0.000 1353.690 4.000 ;
    END
  END lsu_hwdata[55]
  PIN lsu_hwdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 0.000 1359.210 4.000 ;
    END
  END lsu_hwdata[56]
  PIN lsu_hwdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 0.000 1364.270 4.000 ;
    END
  END lsu_hwdata[57]
  PIN lsu_hwdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.510 0.000 1369.790 4.000 ;
    END
  END lsu_hwdata[58]
  PIN lsu_hwdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 0.000 1375.310 4.000 ;
    END
  END lsu_hwdata[59]
  PIN lsu_hwdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 0.000 1083.210 4.000 ;
    END
  END lsu_hwdata[5]
  PIN lsu_hwdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.550 0.000 1380.830 4.000 ;
    END
  END lsu_hwdata[60]
  PIN lsu_hwdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.610 0.000 1385.890 4.000 ;
    END
  END lsu_hwdata[61]
  PIN lsu_hwdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END lsu_hwdata[62]
  PIN lsu_hwdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.650 0.000 1396.930 4.000 ;
    END
  END lsu_hwdata[63]
  PIN lsu_hwdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 0.000 1088.730 4.000 ;
    END
  END lsu_hwdata[6]
  PIN lsu_hwdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.970 0.000 1094.250 4.000 ;
    END
  END lsu_hwdata[7]
  PIN lsu_hwdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.490 0.000 1099.770 4.000 ;
    END
  END lsu_hwdata[8]
  PIN lsu_hwdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END lsu_hwdata[9]
  PIN lsu_hwrite
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END lsu_hwrite
  PIN mbist_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1313.120 4.000 1313.720 ;
    END
  END mbist_mode
  PIN mpc_debug_halt_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1294.760 4.000 1295.360 ;
    END
  END mpc_debug_halt_ack
  PIN mpc_debug_halt_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1290.000 4.000 1290.600 ;
    END
  END mpc_debug_halt_req
  PIN mpc_debug_run_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1296.800 4.000 1297.400 ;
    END
  END mpc_debug_run_ack
  PIN mpc_debug_run_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1291.360 4.000 1291.960 ;
    END
  END mpc_debug_run_req
  PIN mpc_reset_run_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 4.000 1294.000 ;
    END
  END mpc_reset_run_req
  PIN nmi_int
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END nmi_int
  PIN nmi_vec[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END nmi_vec[0]
  PIN nmi_vec[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END nmi_vec[10]
  PIN nmi_vec[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END nmi_vec[11]
  PIN nmi_vec[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END nmi_vec[12]
  PIN nmi_vec[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END nmi_vec[13]
  PIN nmi_vec[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END nmi_vec[14]
  PIN nmi_vec[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END nmi_vec[15]
  PIN nmi_vec[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END nmi_vec[16]
  PIN nmi_vec[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END nmi_vec[17]
  PIN nmi_vec[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END nmi_vec[18]
  PIN nmi_vec[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END nmi_vec[19]
  PIN nmi_vec[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END nmi_vec[1]
  PIN nmi_vec[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END nmi_vec[20]
  PIN nmi_vec[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END nmi_vec[21]
  PIN nmi_vec[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END nmi_vec[22]
  PIN nmi_vec[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END nmi_vec[23]
  PIN nmi_vec[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END nmi_vec[24]
  PIN nmi_vec[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END nmi_vec[25]
  PIN nmi_vec[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END nmi_vec[26]
  PIN nmi_vec[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END nmi_vec[27]
  PIN nmi_vec[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END nmi_vec[28]
  PIN nmi_vec[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END nmi_vec[29]
  PIN nmi_vec[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END nmi_vec[2]
  PIN nmi_vec[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END nmi_vec[30]
  PIN nmi_vec[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END nmi_vec[3]
  PIN nmi_vec[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END nmi_vec[4]
  PIN nmi_vec[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END nmi_vec[5]
  PIN nmi_vec[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END nmi_vec[6]
  PIN nmi_vec[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END nmi_vec[7]
  PIN nmi_vec[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END nmi_vec[8]
  PIN nmi_vec[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END nmi_vec[9]
  PIN o_cpu_halt_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.240 4.000 1302.840 ;
    END
  END o_cpu_halt_ack
  PIN o_cpu_halt_status
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1304.280 4.000 1304.880 ;
    END
  END o_cpu_halt_status
  PIN o_cpu_run_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.040 4.000 1309.640 ;
    END
  END o_cpu_run_ack
  PIN o_debug_mode_status
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1305.640 4.000 1306.240 ;
    END
  END o_debug_mode_status
  PIN rst_l
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END rst_l
  PIN rst_vec[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END rst_vec[0]
  PIN rst_vec[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END rst_vec[10]
  PIN rst_vec[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END rst_vec[11]
  PIN rst_vec[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END rst_vec[12]
  PIN rst_vec[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END rst_vec[13]
  PIN rst_vec[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END rst_vec[14]
  PIN rst_vec[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END rst_vec[15]
  PIN rst_vec[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END rst_vec[16]
  PIN rst_vec[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END rst_vec[17]
  PIN rst_vec[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END rst_vec[18]
  PIN rst_vec[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END rst_vec[19]
  PIN rst_vec[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END rst_vec[1]
  PIN rst_vec[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END rst_vec[20]
  PIN rst_vec[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END rst_vec[21]
  PIN rst_vec[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END rst_vec[22]
  PIN rst_vec[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END rst_vec[23]
  PIN rst_vec[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END rst_vec[24]
  PIN rst_vec[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END rst_vec[25]
  PIN rst_vec[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END rst_vec[26]
  PIN rst_vec[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END rst_vec[27]
  PIN rst_vec[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END rst_vec[28]
  PIN rst_vec[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END rst_vec[29]
  PIN rst_vec[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END rst_vec[2]
  PIN rst_vec[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END rst_vec[30]
  PIN rst_vec[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END rst_vec[3]
  PIN rst_vec[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END rst_vec[4]
  PIN rst_vec[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END rst_vec[5]
  PIN rst_vec[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END rst_vec[6]
  PIN rst_vec[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END rst_vec[7]
  PIN rst_vec[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END rst_vec[8]
  PIN rst_vec[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END rst_vec[9]
  PIN sb_haddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END sb_haddr[0]
  PIN sb_haddr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.880 4.000 247.480 ;
    END
  END sb_haddr[10]
  PIN sb_haddr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END sb_haddr[11]
  PIN sb_haddr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END sb_haddr[12]
  PIN sb_haddr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END sb_haddr[13]
  PIN sb_haddr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END sb_haddr[14]
  PIN sb_haddr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END sb_haddr[15]
  PIN sb_haddr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END sb_haddr[16]
  PIN sb_haddr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END sb_haddr[17]
  PIN sb_haddr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END sb_haddr[18]
  PIN sb_haddr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END sb_haddr[19]
  PIN sb_haddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END sb_haddr[1]
  PIN sb_haddr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END sb_haddr[20]
  PIN sb_haddr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END sb_haddr[21]
  PIN sb_haddr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END sb_haddr[22]
  PIN sb_haddr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END sb_haddr[23]
  PIN sb_haddr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END sb_haddr[24]
  PIN sb_haddr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END sb_haddr[25]
  PIN sb_haddr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END sb_haddr[26]
  PIN sb_haddr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END sb_haddr[27]
  PIN sb_haddr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END sb_haddr[28]
  PIN sb_haddr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END sb_haddr[29]
  PIN sb_haddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END sb_haddr[2]
  PIN sb_haddr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END sb_haddr[30]
  PIN sb_haddr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END sb_haddr[31]
  PIN sb_haddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END sb_haddr[3]
  PIN sb_haddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END sb_haddr[4]
  PIN sb_haddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END sb_haddr[5]
  PIN sb_haddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END sb_haddr[6]
  PIN sb_haddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END sb_haddr[7]
  PIN sb_haddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END sb_haddr[8]
  PIN sb_haddr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END sb_haddr[9]
  PIN sb_hburst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END sb_hburst[0]
  PIN sb_hburst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END sb_hburst[1]
  PIN sb_hburst[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END sb_hburst[2]
  PIN sb_hmastlock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END sb_hmastlock
  PIN sb_hprot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END sb_hprot[0]
  PIN sb_hprot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END sb_hprot[1]
  PIN sb_hprot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END sb_hprot[2]
  PIN sb_hprot[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END sb_hprot[3]
  PIN sb_hrdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END sb_hrdata[0]
  PIN sb_hrdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END sb_hrdata[10]
  PIN sb_hrdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END sb_hrdata[11]
  PIN sb_hrdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.800 4.000 447.400 ;
    END
  END sb_hrdata[12]
  PIN sb_hrdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END sb_hrdata[13]
  PIN sb_hrdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END sb_hrdata[14]
  PIN sb_hrdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END sb_hrdata[15]
  PIN sb_hrdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END sb_hrdata[16]
  PIN sb_hrdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END sb_hrdata[17]
  PIN sb_hrdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END sb_hrdata[18]
  PIN sb_hrdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END sb_hrdata[19]
  PIN sb_hrdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END sb_hrdata[1]
  PIN sb_hrdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END sb_hrdata[20]
  PIN sb_hrdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END sb_hrdata[21]
  PIN sb_hrdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 464.480 4.000 465.080 ;
    END
  END sb_hrdata[22]
  PIN sb_hrdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END sb_hrdata[23]
  PIN sb_hrdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END sb_hrdata[24]
  PIN sb_hrdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.920 4.000 470.520 ;
    END
  END sb_hrdata[25]
  PIN sb_hrdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END sb_hrdata[26]
  PIN sb_hrdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END sb_hrdata[27]
  PIN sb_hrdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 475.360 4.000 475.960 ;
    END
  END sb_hrdata[28]
  PIN sb_hrdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END sb_hrdata[29]
  PIN sb_hrdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END sb_hrdata[2]
  PIN sb_hrdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END sb_hrdata[30]
  PIN sb_hrdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END sb_hrdata[31]
  PIN sb_hrdata[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END sb_hrdata[32]
  PIN sb_hrdata[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END sb_hrdata[33]
  PIN sb_hrdata[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END sb_hrdata[34]
  PIN sb_hrdata[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 487.600 4.000 488.200 ;
    END
  END sb_hrdata[35]
  PIN sb_hrdata[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END sb_hrdata[36]
  PIN sb_hrdata[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.680 4.000 492.280 ;
    END
  END sb_hrdata[37]
  PIN sb_hrdata[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END sb_hrdata[38]
  PIN sb_hrdata[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END sb_hrdata[39]
  PIN sb_hrdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END sb_hrdata[3]
  PIN sb_hrdata[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.120 4.000 497.720 ;
    END
  END sb_hrdata[40]
  PIN sb_hrdata[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 498.480 4.000 499.080 ;
    END
  END sb_hrdata[41]
  PIN sb_hrdata[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END sb_hrdata[42]
  PIN sb_hrdata[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END sb_hrdata[43]
  PIN sb_hrdata[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.920 4.000 504.520 ;
    END
  END sb_hrdata[44]
  PIN sb_hrdata[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END sb_hrdata[45]
  PIN sb_hrdata[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END sb_hrdata[46]
  PIN sb_hrdata[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 509.360 4.000 509.960 ;
    END
  END sb_hrdata[47]
  PIN sb_hrdata[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END sb_hrdata[48]
  PIN sb_hrdata[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END sb_hrdata[49]
  PIN sb_hrdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END sb_hrdata[4]
  PIN sb_hrdata[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END sb_hrdata[50]
  PIN sb_hrdata[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.160 4.000 516.760 ;
    END
  END sb_hrdata[51]
  PIN sb_hrdata[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END sb_hrdata[52]
  PIN sb_hrdata[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END sb_hrdata[53]
  PIN sb_hrdata[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 521.600 4.000 522.200 ;
    END
  END sb_hrdata[54]
  PIN sb_hrdata[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END sb_hrdata[55]
  PIN sb_hrdata[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.680 4.000 526.280 ;
    END
  END sb_hrdata[56]
  PIN sb_hrdata[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END sb_hrdata[57]
  PIN sb_hrdata[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END sb_hrdata[58]
  PIN sb_hrdata[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END sb_hrdata[59]
  PIN sb_hrdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.560 4.000 435.160 ;
    END
  END sb_hrdata[5]
  PIN sb_hrdata[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 532.480 4.000 533.080 ;
    END
  END sb_hrdata[60]
  PIN sb_hrdata[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END sb_hrdata[61]
  PIN sb_hrdata[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END sb_hrdata[62]
  PIN sb_hrdata[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.920 4.000 538.520 ;
    END
  END sb_hrdata[63]
  PIN sb_hrdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.920 4.000 436.520 ;
    END
  END sb_hrdata[6]
  PIN sb_hrdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END sb_hrdata[7]
  PIN sb_hrdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END sb_hrdata[8]
  PIN sb_hrdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END sb_hrdata[9]
  PIN sb_hready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END sb_hready
  PIN sb_hresp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END sb_hresp
  PIN sb_hsize[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END sb_hsize[0]
  PIN sb_hsize[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END sb_hsize[1]
  PIN sb_hsize[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END sb_hsize[2]
  PIN sb_htrans[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END sb_htrans[0]
  PIN sb_htrans[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END sb_htrans[1]
  PIN sb_hwdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END sb_hwdata[0]
  PIN sb_hwdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END sb_hwdata[10]
  PIN sb_hwdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END sb_hwdata[11]
  PIN sb_hwdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.560 4.000 333.160 ;
    END
  END sb_hwdata[12]
  PIN sb_hwdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END sb_hwdata[13]
  PIN sb_hwdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END sb_hwdata[14]
  PIN sb_hwdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END sb_hwdata[15]
  PIN sb_hwdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END sb_hwdata[16]
  PIN sb_hwdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END sb_hwdata[17]
  PIN sb_hwdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END sb_hwdata[18]
  PIN sb_hwdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END sb_hwdata[19]
  PIN sb_hwdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END sb_hwdata[1]
  PIN sb_hwdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END sb_hwdata[20]
  PIN sb_hwdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END sb_hwdata[21]
  PIN sb_hwdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END sb_hwdata[22]
  PIN sb_hwdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END sb_hwdata[23]
  PIN sb_hwdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END sb_hwdata[24]
  PIN sb_hwdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END sb_hwdata[25]
  PIN sb_hwdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END sb_hwdata[26]
  PIN sb_hwdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END sb_hwdata[27]
  PIN sb_hwdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END sb_hwdata[28]
  PIN sb_hwdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END sb_hwdata[29]
  PIN sb_hwdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END sb_hwdata[2]
  PIN sb_hwdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END sb_hwdata[30]
  PIN sb_hwdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END sb_hwdata[31]
  PIN sb_hwdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END sb_hwdata[32]
  PIN sb_hwdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END sb_hwdata[33]
  PIN sb_hwdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.000 4.000 372.600 ;
    END
  END sb_hwdata[34]
  PIN sb_hwdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END sb_hwdata[35]
  PIN sb_hwdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END sb_hwdata[36]
  PIN sb_hwdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END sb_hwdata[37]
  PIN sb_hwdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END sb_hwdata[38]
  PIN sb_hwdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END sb_hwdata[39]
  PIN sb_hwdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END sb_hwdata[3]
  PIN sb_hwdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END sb_hwdata[40]
  PIN sb_hwdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END sb_hwdata[41]
  PIN sb_hwdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END sb_hwdata[42]
  PIN sb_hwdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END sb_hwdata[43]
  PIN sb_hwdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END sb_hwdata[44]
  PIN sb_hwdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END sb_hwdata[45]
  PIN sb_hwdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END sb_hwdata[46]
  PIN sb_hwdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END sb_hwdata[47]
  PIN sb_hwdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END sb_hwdata[48]
  PIN sb_hwdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END sb_hwdata[49]
  PIN sb_hwdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END sb_hwdata[4]
  PIN sb_hwdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.560 4.000 401.160 ;
    END
  END sb_hwdata[50]
  PIN sb_hwdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END sb_hwdata[51]
  PIN sb_hwdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END sb_hwdata[52]
  PIN sb_hwdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END sb_hwdata[53]
  PIN sb_hwdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END sb_hwdata[54]
  PIN sb_hwdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END sb_hwdata[55]
  PIN sb_hwdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END sb_hwdata[56]
  PIN sb_hwdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END sb_hwdata[57]
  PIN sb_hwdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END sb_hwdata[58]
  PIN sb_hwdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END sb_hwdata[59]
  PIN sb_hwdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END sb_hwdata[5]
  PIN sb_hwdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END sb_hwdata[60]
  PIN sb_hwdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END sb_hwdata[61]
  PIN sb_hwdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END sb_hwdata[62]
  PIN sb_hwdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END sb_hwdata[63]
  PIN sb_hwdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END sb_hwdata[6]
  PIN sb_hwdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END sb_hwdata[7]
  PIN sb_hwdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END sb_hwdata[8]
  PIN sb_hwdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END sb_hwdata[9]
  PIN sb_hwrite
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END sb_hwrite
  PIN scan_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1311.080 4.000 1311.680 ;
    END
  END scan_mode
  PIN soft_int
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END soft_int
  PIN timer_int
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END timer_int
  PIN trace_rv_i_address_ip[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1314.480 4.000 1315.080 ;
    END
  END trace_rv_i_address_ip[0]
  PIN trace_rv_i_address_ip[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END trace_rv_i_address_ip[10]
  PIN trace_rv_i_address_ip[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1334.200 4.000 1334.800 ;
    END
  END trace_rv_i_address_ip[11]
  PIN trace_rv_i_address_ip[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1336.240 4.000 1336.840 ;
    END
  END trace_rv_i_address_ip[12]
  PIN trace_rv_i_address_ip[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1338.280 4.000 1338.880 ;
    END
  END trace_rv_i_address_ip[13]
  PIN trace_rv_i_address_ip[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1339.640 4.000 1340.240 ;
    END
  END trace_rv_i_address_ip[14]
  PIN trace_rv_i_address_ip[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1341.680 4.000 1342.280 ;
    END
  END trace_rv_i_address_ip[15]
  PIN trace_rv_i_address_ip[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.040 4.000 1343.640 ;
    END
  END trace_rv_i_address_ip[16]
  PIN trace_rv_i_address_ip[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1345.080 4.000 1345.680 ;
    END
  END trace_rv_i_address_ip[17]
  PIN trace_rv_i_address_ip[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1347.120 4.000 1347.720 ;
    END
  END trace_rv_i_address_ip[18]
  PIN trace_rv_i_address_ip[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1348.480 4.000 1349.080 ;
    END
  END trace_rv_i_address_ip[19]
  PIN trace_rv_i_address_ip[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1316.520 4.000 1317.120 ;
    END
  END trace_rv_i_address_ip[1]
  PIN trace_rv_i_address_ip[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1350.520 4.000 1351.120 ;
    END
  END trace_rv_i_address_ip[20]
  PIN trace_rv_i_address_ip[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1352.560 4.000 1353.160 ;
    END
  END trace_rv_i_address_ip[21]
  PIN trace_rv_i_address_ip[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.920 4.000 1354.520 ;
    END
  END trace_rv_i_address_ip[22]
  PIN trace_rv_i_address_ip[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1355.960 4.000 1356.560 ;
    END
  END trace_rv_i_address_ip[23]
  PIN trace_rv_i_address_ip[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1357.320 4.000 1357.920 ;
    END
  END trace_rv_i_address_ip[24]
  PIN trace_rv_i_address_ip[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1359.360 4.000 1359.960 ;
    END
  END trace_rv_i_address_ip[25]
  PIN trace_rv_i_address_ip[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1361.400 4.000 1362.000 ;
    END
  END trace_rv_i_address_ip[26]
  PIN trace_rv_i_address_ip[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1362.760 4.000 1363.360 ;
    END
  END trace_rv_i_address_ip[27]
  PIN trace_rv_i_address_ip[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1364.800 4.000 1365.400 ;
    END
  END trace_rv_i_address_ip[28]
  PIN trace_rv_i_address_ip[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1366.840 4.000 1367.440 ;
    END
  END trace_rv_i_address_ip[29]
  PIN trace_rv_i_address_ip[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1318.560 4.000 1319.160 ;
    END
  END trace_rv_i_address_ip[2]
  PIN trace_rv_i_address_ip[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1368.200 4.000 1368.800 ;
    END
  END trace_rv_i_address_ip[30]
  PIN trace_rv_i_address_ip[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.240 4.000 1370.840 ;
    END
  END trace_rv_i_address_ip[31]
  PIN trace_rv_i_address_ip[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1319.920 4.000 1320.520 ;
    END
  END trace_rv_i_address_ip[3]
  PIN trace_rv_i_address_ip[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1321.960 4.000 1322.560 ;
    END
  END trace_rv_i_address_ip[4]
  PIN trace_rv_i_address_ip[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1324.000 4.000 1324.600 ;
    END
  END trace_rv_i_address_ip[5]
  PIN trace_rv_i_address_ip[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1325.360 4.000 1325.960 ;
    END
  END trace_rv_i_address_ip[6]
  PIN trace_rv_i_address_ip[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1327.400 4.000 1328.000 ;
    END
  END trace_rv_i_address_ip[7]
  PIN trace_rv_i_address_ip[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1328.760 4.000 1329.360 ;
    END
  END trace_rv_i_address_ip[8]
  PIN trace_rv_i_address_ip[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1330.800 4.000 1331.400 ;
    END
  END trace_rv_i_address_ip[9]
  PIN trace_rv_i_ecause_ip[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1371.600 4.000 1372.200 ;
    END
  END trace_rv_i_ecause_ip[0]
  PIN trace_rv_i_ecause_ip[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1373.640 4.000 1374.240 ;
    END
  END trace_rv_i_ecause_ip[1]
  PIN trace_rv_i_ecause_ip[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1375.680 4.000 1376.280 ;
    END
  END trace_rv_i_ecause_ip[2]
  PIN trace_rv_i_ecause_ip[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.040 4.000 1377.640 ;
    END
  END trace_rv_i_ecause_ip[3]
  PIN trace_rv_i_ecause_ip[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1379.080 4.000 1379.680 ;
    END
  END trace_rv_i_ecause_ip[4]
  PIN trace_rv_i_exception_ip
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1381.120 4.000 1381.720 ;
    END
  END trace_rv_i_exception_ip
  PIN trace_rv_i_insn_ip[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1382.480 4.000 1383.080 ;
    END
  END trace_rv_i_insn_ip[0]
  PIN trace_rv_i_insn_ip[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1400.160 4.000 1400.760 ;
    END
  END trace_rv_i_insn_ip[10]
  PIN trace_rv_i_insn_ip[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1402.200 4.000 1402.800 ;
    END
  END trace_rv_i_insn_ip[11]
  PIN trace_rv_i_insn_ip[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1404.240 4.000 1404.840 ;
    END
  END trace_rv_i_insn_ip[12]
  PIN trace_rv_i_insn_ip[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1405.600 4.000 1406.200 ;
    END
  END trace_rv_i_insn_ip[13]
  PIN trace_rv_i_insn_ip[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 4.000 1408.240 ;
    END
  END trace_rv_i_insn_ip[14]
  PIN trace_rv_i_insn_ip[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1409.680 4.000 1410.280 ;
    END
  END trace_rv_i_insn_ip[15]
  PIN trace_rv_i_insn_ip[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.040 4.000 1411.640 ;
    END
  END trace_rv_i_insn_ip[16]
  PIN trace_rv_i_insn_ip[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1413.080 4.000 1413.680 ;
    END
  END trace_rv_i_insn_ip[17]
  PIN trace_rv_i_insn_ip[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1414.440 4.000 1415.040 ;
    END
  END trace_rv_i_insn_ip[18]
  PIN trace_rv_i_insn_ip[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1416.480 4.000 1417.080 ;
    END
  END trace_rv_i_insn_ip[19]
  PIN trace_rv_i_insn_ip[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1384.520 4.000 1385.120 ;
    END
  END trace_rv_i_insn_ip[1]
  PIN trace_rv_i_insn_ip[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1418.520 4.000 1419.120 ;
    END
  END trace_rv_i_insn_ip[20]
  PIN trace_rv_i_insn_ip[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1419.880 4.000 1420.480 ;
    END
  END trace_rv_i_insn_ip[21]
  PIN trace_rv_i_insn_ip[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1421.920 4.000 1422.520 ;
    END
  END trace_rv_i_insn_ip[22]
  PIN trace_rv_i_insn_ip[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1423.960 4.000 1424.560 ;
    END
  END trace_rv_i_insn_ip[23]
  PIN trace_rv_i_insn_ip[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1425.320 4.000 1425.920 ;
    END
  END trace_rv_i_insn_ip[24]
  PIN trace_rv_i_insn_ip[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1427.360 4.000 1427.960 ;
    END
  END trace_rv_i_insn_ip[25]
  PIN trace_rv_i_insn_ip[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1428.720 4.000 1429.320 ;
    END
  END trace_rv_i_insn_ip[26]
  PIN trace_rv_i_insn_ip[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1430.760 4.000 1431.360 ;
    END
  END trace_rv_i_insn_ip[27]
  PIN trace_rv_i_insn_ip[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1432.800 4.000 1433.400 ;
    END
  END trace_rv_i_insn_ip[28]
  PIN trace_rv_i_insn_ip[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.160 4.000 1434.760 ;
    END
  END trace_rv_i_insn_ip[29]
  PIN trace_rv_i_insn_ip[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1385.880 4.000 1386.480 ;
    END
  END trace_rv_i_insn_ip[2]
  PIN trace_rv_i_insn_ip[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1436.200 4.000 1436.800 ;
    END
  END trace_rv_i_insn_ip[30]
  PIN trace_rv_i_insn_ip[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1438.240 4.000 1438.840 ;
    END
  END trace_rv_i_insn_ip[31]
  PIN trace_rv_i_insn_ip[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1387.920 4.000 1388.520 ;
    END
  END trace_rv_i_insn_ip[3]
  PIN trace_rv_i_insn_ip[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1389.960 4.000 1390.560 ;
    END
  END trace_rv_i_insn_ip[4]
  PIN trace_rv_i_insn_ip[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1391.320 4.000 1391.920 ;
    END
  END trace_rv_i_insn_ip[5]
  PIN trace_rv_i_insn_ip[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1393.360 4.000 1393.960 ;
    END
  END trace_rv_i_insn_ip[6]
  PIN trace_rv_i_insn_ip[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1395.400 4.000 1396.000 ;
    END
  END trace_rv_i_insn_ip[7]
  PIN trace_rv_i_insn_ip[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1396.760 4.000 1397.360 ;
    END
  END trace_rv_i_insn_ip[8]
  PIN trace_rv_i_insn_ip[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1398.800 4.000 1399.400 ;
    END
  END trace_rv_i_insn_ip[9]
  PIN trace_rv_i_interrupt_ip
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1439.600 4.000 1440.200 ;
    END
  END trace_rv_i_interrupt_ip
  PIN trace_rv_i_tval_ip[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1441.640 4.000 1442.240 ;
    END
  END trace_rv_i_tval_ip[0]
  PIN trace_rv_i_tval_ip[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1459.320 4.000 1459.920 ;
    END
  END trace_rv_i_tval_ip[10]
  PIN trace_rv_i_tval_ip[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1461.360 4.000 1461.960 ;
    END
  END trace_rv_i_tval_ip[11]
  PIN trace_rv_i_tval_ip[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.720 4.000 1463.320 ;
    END
  END trace_rv_i_tval_ip[12]
  PIN trace_rv_i_tval_ip[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1464.760 4.000 1465.360 ;
    END
  END trace_rv_i_tval_ip[13]
  PIN trace_rv_i_tval_ip[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1466.800 4.000 1467.400 ;
    END
  END trace_rv_i_tval_ip[14]
  PIN trace_rv_i_tval_ip[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1468.160 4.000 1468.760 ;
    END
  END trace_rv_i_tval_ip[15]
  PIN trace_rv_i_tval_ip[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1470.200 4.000 1470.800 ;
    END
  END trace_rv_i_tval_ip[16]
  PIN trace_rv_i_tval_ip[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1471.560 4.000 1472.160 ;
    END
  END trace_rv_i_tval_ip[17]
  PIN trace_rv_i_tval_ip[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1473.600 4.000 1474.200 ;
    END
  END trace_rv_i_tval_ip[18]
  PIN trace_rv_i_tval_ip[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1475.640 4.000 1476.240 ;
    END
  END trace_rv_i_tval_ip[19]
  PIN trace_rv_i_tval_ip[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1443.000 4.000 1443.600 ;
    END
  END trace_rv_i_tval_ip[1]
  PIN trace_rv_i_tval_ip[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1477.000 4.000 1477.600 ;
    END
  END trace_rv_i_tval_ip[20]
  PIN trace_rv_i_tval_ip[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1479.040 4.000 1479.640 ;
    END
  END trace_rv_i_tval_ip[21]
  PIN trace_rv_i_tval_ip[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1481.080 4.000 1481.680 ;
    END
  END trace_rv_i_tval_ip[22]
  PIN trace_rv_i_tval_ip[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1482.440 4.000 1483.040 ;
    END
  END trace_rv_i_tval_ip[23]
  PIN trace_rv_i_tval_ip[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1484.480 4.000 1485.080 ;
    END
  END trace_rv_i_tval_ip[24]
  PIN trace_rv_i_tval_ip[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1485.840 4.000 1486.440 ;
    END
  END trace_rv_i_tval_ip[25]
  PIN trace_rv_i_tval_ip[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1487.880 4.000 1488.480 ;
    END
  END trace_rv_i_tval_ip[26]
  PIN trace_rv_i_tval_ip[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.920 4.000 1490.520 ;
    END
  END trace_rv_i_tval_ip[27]
  PIN trace_rv_i_tval_ip[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1491.280 4.000 1491.880 ;
    END
  END trace_rv_i_tval_ip[28]
  PIN trace_rv_i_tval_ip[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1493.320 4.000 1493.920 ;
    END
  END trace_rv_i_tval_ip[29]
  PIN trace_rv_i_tval_ip[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.040 4.000 1445.640 ;
    END
  END trace_rv_i_tval_ip[2]
  PIN trace_rv_i_tval_ip[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1495.360 4.000 1495.960 ;
    END
  END trace_rv_i_tval_ip[30]
  PIN trace_rv_i_tval_ip[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1496.720 4.000 1497.320 ;
    END
  END trace_rv_i_tval_ip[31]
  PIN trace_rv_i_tval_ip[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1447.080 4.000 1447.680 ;
    END
  END trace_rv_i_tval_ip[3]
  PIN trace_rv_i_tval_ip[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1448.440 4.000 1449.040 ;
    END
  END trace_rv_i_tval_ip[4]
  PIN trace_rv_i_tval_ip[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1450.480 4.000 1451.080 ;
    END
  END trace_rv_i_tval_ip[5]
  PIN trace_rv_i_tval_ip[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1452.520 4.000 1453.120 ;
    END
  END trace_rv_i_tval_ip[6]
  PIN trace_rv_i_tval_ip[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1453.880 4.000 1454.480 ;
    END
  END trace_rv_i_tval_ip[7]
  PIN trace_rv_i_tval_ip[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.920 4.000 1456.520 ;
    END
  END trace_rv_i_tval_ip[8]
  PIN trace_rv_i_tval_ip[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1457.280 4.000 1457.880 ;
    END
  END trace_rv_i_tval_ip[9]
  PIN trace_rv_i_valid_ip
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1498.760 4.000 1499.360 ;
    END
  END trace_rv_i_valid_ip
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.745 10.795 1394.260 1487.925 ;
      LAYER met1 ;
        RECT 0.070 0.040 1396.950 1490.860 ;
      LAYER met2 ;
        RECT 0.100 4.280 1396.920 1499.245 ;
        RECT 0.100 0.010 2.110 4.280 ;
        RECT 2.950 0.010 7.170 4.280 ;
        RECT 8.010 0.010 12.690 4.280 ;
        RECT 13.530 0.010 18.210 4.280 ;
        RECT 19.050 0.010 23.270 4.280 ;
        RECT 24.110 0.010 28.790 4.280 ;
        RECT 29.630 0.010 34.310 4.280 ;
        RECT 35.150 0.010 39.830 4.280 ;
        RECT 40.670 0.010 44.890 4.280 ;
        RECT 45.730 0.010 50.410 4.280 ;
        RECT 51.250 0.010 55.930 4.280 ;
        RECT 56.770 0.010 61.450 4.280 ;
        RECT 62.290 0.010 66.510 4.280 ;
        RECT 67.350 0.010 72.030 4.280 ;
        RECT 72.870 0.010 77.550 4.280 ;
        RECT 78.390 0.010 83.070 4.280 ;
        RECT 83.910 0.010 88.130 4.280 ;
        RECT 88.970 0.010 93.650 4.280 ;
        RECT 94.490 0.010 99.170 4.280 ;
        RECT 100.010 0.010 104.690 4.280 ;
        RECT 105.530 0.010 109.750 4.280 ;
        RECT 110.590 0.010 115.270 4.280 ;
        RECT 116.110 0.010 120.790 4.280 ;
        RECT 121.630 0.010 126.310 4.280 ;
        RECT 127.150 0.010 131.370 4.280 ;
        RECT 132.210 0.010 136.890 4.280 ;
        RECT 137.730 0.010 142.410 4.280 ;
        RECT 143.250 0.010 147.930 4.280 ;
        RECT 148.770 0.010 152.990 4.280 ;
        RECT 153.830 0.010 158.510 4.280 ;
        RECT 159.350 0.010 164.030 4.280 ;
        RECT 164.870 0.010 169.550 4.280 ;
        RECT 170.390 0.010 174.610 4.280 ;
        RECT 175.450 0.010 180.130 4.280 ;
        RECT 180.970 0.010 185.650 4.280 ;
        RECT 186.490 0.010 191.170 4.280 ;
        RECT 192.010 0.010 196.230 4.280 ;
        RECT 197.070 0.010 201.750 4.280 ;
        RECT 202.590 0.010 207.270 4.280 ;
        RECT 208.110 0.010 212.790 4.280 ;
        RECT 213.630 0.010 217.850 4.280 ;
        RECT 218.690 0.010 223.370 4.280 ;
        RECT 224.210 0.010 228.890 4.280 ;
        RECT 229.730 0.010 234.410 4.280 ;
        RECT 235.250 0.010 239.470 4.280 ;
        RECT 240.310 0.010 244.990 4.280 ;
        RECT 245.830 0.010 250.510 4.280 ;
        RECT 251.350 0.010 256.030 4.280 ;
        RECT 256.870 0.010 261.090 4.280 ;
        RECT 261.930 0.010 266.610 4.280 ;
        RECT 267.450 0.010 272.130 4.280 ;
        RECT 272.970 0.010 277.650 4.280 ;
        RECT 278.490 0.010 282.710 4.280 ;
        RECT 283.550 0.010 288.230 4.280 ;
        RECT 289.070 0.010 293.750 4.280 ;
        RECT 294.590 0.010 299.270 4.280 ;
        RECT 300.110 0.010 304.330 4.280 ;
        RECT 305.170 0.010 309.850 4.280 ;
        RECT 310.690 0.010 315.370 4.280 ;
        RECT 316.210 0.010 320.890 4.280 ;
        RECT 321.730 0.010 325.950 4.280 ;
        RECT 326.790 0.010 331.470 4.280 ;
        RECT 332.310 0.010 336.990 4.280 ;
        RECT 337.830 0.010 342.510 4.280 ;
        RECT 343.350 0.010 347.570 4.280 ;
        RECT 348.410 0.010 353.090 4.280 ;
        RECT 353.930 0.010 358.610 4.280 ;
        RECT 359.450 0.010 364.130 4.280 ;
        RECT 364.970 0.010 369.190 4.280 ;
        RECT 370.030 0.010 374.710 4.280 ;
        RECT 375.550 0.010 380.230 4.280 ;
        RECT 381.070 0.010 385.750 4.280 ;
        RECT 386.590 0.010 390.810 4.280 ;
        RECT 391.650 0.010 396.330 4.280 ;
        RECT 397.170 0.010 401.850 4.280 ;
        RECT 402.690 0.010 407.370 4.280 ;
        RECT 408.210 0.010 412.430 4.280 ;
        RECT 413.270 0.010 417.950 4.280 ;
        RECT 418.790 0.010 423.470 4.280 ;
        RECT 424.310 0.010 428.990 4.280 ;
        RECT 429.830 0.010 434.050 4.280 ;
        RECT 434.890 0.010 439.570 4.280 ;
        RECT 440.410 0.010 445.090 4.280 ;
        RECT 445.930 0.010 450.610 4.280 ;
        RECT 451.450 0.010 455.670 4.280 ;
        RECT 456.510 0.010 461.190 4.280 ;
        RECT 462.030 0.010 466.710 4.280 ;
        RECT 467.550 0.010 472.230 4.280 ;
        RECT 473.070 0.010 477.290 4.280 ;
        RECT 478.130 0.010 482.810 4.280 ;
        RECT 483.650 0.010 488.330 4.280 ;
        RECT 489.170 0.010 493.850 4.280 ;
        RECT 494.690 0.010 498.910 4.280 ;
        RECT 499.750 0.010 504.430 4.280 ;
        RECT 505.270 0.010 509.950 4.280 ;
        RECT 510.790 0.010 515.470 4.280 ;
        RECT 516.310 0.010 520.530 4.280 ;
        RECT 521.370 0.010 526.050 4.280 ;
        RECT 526.890 0.010 531.570 4.280 ;
        RECT 532.410 0.010 537.090 4.280 ;
        RECT 537.930 0.010 542.150 4.280 ;
        RECT 542.990 0.010 547.670 4.280 ;
        RECT 548.510 0.010 553.190 4.280 ;
        RECT 554.030 0.010 558.710 4.280 ;
        RECT 559.550 0.010 563.770 4.280 ;
        RECT 564.610 0.010 569.290 4.280 ;
        RECT 570.130 0.010 574.810 4.280 ;
        RECT 575.650 0.010 580.330 4.280 ;
        RECT 581.170 0.010 585.390 4.280 ;
        RECT 586.230 0.010 590.910 4.280 ;
        RECT 591.750 0.010 596.430 4.280 ;
        RECT 597.270 0.010 601.950 4.280 ;
        RECT 602.790 0.010 607.010 4.280 ;
        RECT 607.850 0.010 612.530 4.280 ;
        RECT 613.370 0.010 618.050 4.280 ;
        RECT 618.890 0.010 623.570 4.280 ;
        RECT 624.410 0.010 628.630 4.280 ;
        RECT 629.470 0.010 634.150 4.280 ;
        RECT 634.990 0.010 639.670 4.280 ;
        RECT 640.510 0.010 645.190 4.280 ;
        RECT 646.030 0.010 650.250 4.280 ;
        RECT 651.090 0.010 655.770 4.280 ;
        RECT 656.610 0.010 661.290 4.280 ;
        RECT 662.130 0.010 666.810 4.280 ;
        RECT 667.650 0.010 671.870 4.280 ;
        RECT 672.710 0.010 677.390 4.280 ;
        RECT 678.230 0.010 682.910 4.280 ;
        RECT 683.750 0.010 688.430 4.280 ;
        RECT 689.270 0.010 693.490 4.280 ;
        RECT 694.330 0.010 699.010 4.280 ;
        RECT 699.850 0.010 704.530 4.280 ;
        RECT 705.370 0.010 710.050 4.280 ;
        RECT 710.890 0.010 715.110 4.280 ;
        RECT 715.950 0.010 720.630 4.280 ;
        RECT 721.470 0.010 726.150 4.280 ;
        RECT 726.990 0.010 731.670 4.280 ;
        RECT 732.510 0.010 736.730 4.280 ;
        RECT 737.570 0.010 742.250 4.280 ;
        RECT 743.090 0.010 747.770 4.280 ;
        RECT 748.610 0.010 753.290 4.280 ;
        RECT 754.130 0.010 758.350 4.280 ;
        RECT 759.190 0.010 763.870 4.280 ;
        RECT 764.710 0.010 769.390 4.280 ;
        RECT 770.230 0.010 774.910 4.280 ;
        RECT 775.750 0.010 779.970 4.280 ;
        RECT 780.810 0.010 785.490 4.280 ;
        RECT 786.330 0.010 791.010 4.280 ;
        RECT 791.850 0.010 796.530 4.280 ;
        RECT 797.370 0.010 801.590 4.280 ;
        RECT 802.430 0.010 807.110 4.280 ;
        RECT 807.950 0.010 812.630 4.280 ;
        RECT 813.470 0.010 818.150 4.280 ;
        RECT 818.990 0.010 823.210 4.280 ;
        RECT 824.050 0.010 828.730 4.280 ;
        RECT 829.570 0.010 834.250 4.280 ;
        RECT 835.090 0.010 839.770 4.280 ;
        RECT 840.610 0.010 844.830 4.280 ;
        RECT 845.670 0.010 850.350 4.280 ;
        RECT 851.190 0.010 855.870 4.280 ;
        RECT 856.710 0.010 861.390 4.280 ;
        RECT 862.230 0.010 866.450 4.280 ;
        RECT 867.290 0.010 871.970 4.280 ;
        RECT 872.810 0.010 877.490 4.280 ;
        RECT 878.330 0.010 883.010 4.280 ;
        RECT 883.850 0.010 888.070 4.280 ;
        RECT 888.910 0.010 893.590 4.280 ;
        RECT 894.430 0.010 899.110 4.280 ;
        RECT 899.950 0.010 904.630 4.280 ;
        RECT 905.470 0.010 909.690 4.280 ;
        RECT 910.530 0.010 915.210 4.280 ;
        RECT 916.050 0.010 920.730 4.280 ;
        RECT 921.570 0.010 926.250 4.280 ;
        RECT 927.090 0.010 931.310 4.280 ;
        RECT 932.150 0.010 936.830 4.280 ;
        RECT 937.670 0.010 942.350 4.280 ;
        RECT 943.190 0.010 947.870 4.280 ;
        RECT 948.710 0.010 952.930 4.280 ;
        RECT 953.770 0.010 958.450 4.280 ;
        RECT 959.290 0.010 963.970 4.280 ;
        RECT 964.810 0.010 969.490 4.280 ;
        RECT 970.330 0.010 974.550 4.280 ;
        RECT 975.390 0.010 980.070 4.280 ;
        RECT 980.910 0.010 985.590 4.280 ;
        RECT 986.430 0.010 991.110 4.280 ;
        RECT 991.950 0.010 996.170 4.280 ;
        RECT 997.010 0.010 1001.690 4.280 ;
        RECT 1002.530 0.010 1007.210 4.280 ;
        RECT 1008.050 0.010 1012.730 4.280 ;
        RECT 1013.570 0.010 1017.790 4.280 ;
        RECT 1018.630 0.010 1023.310 4.280 ;
        RECT 1024.150 0.010 1028.830 4.280 ;
        RECT 1029.670 0.010 1034.350 4.280 ;
        RECT 1035.190 0.010 1039.410 4.280 ;
        RECT 1040.250 0.010 1044.930 4.280 ;
        RECT 1045.770 0.010 1050.450 4.280 ;
        RECT 1051.290 0.010 1055.970 4.280 ;
        RECT 1056.810 0.010 1061.030 4.280 ;
        RECT 1061.870 0.010 1066.550 4.280 ;
        RECT 1067.390 0.010 1072.070 4.280 ;
        RECT 1072.910 0.010 1077.590 4.280 ;
        RECT 1078.430 0.010 1082.650 4.280 ;
        RECT 1083.490 0.010 1088.170 4.280 ;
        RECT 1089.010 0.010 1093.690 4.280 ;
        RECT 1094.530 0.010 1099.210 4.280 ;
        RECT 1100.050 0.010 1104.270 4.280 ;
        RECT 1105.110 0.010 1109.790 4.280 ;
        RECT 1110.630 0.010 1115.310 4.280 ;
        RECT 1116.150 0.010 1120.830 4.280 ;
        RECT 1121.670 0.010 1125.890 4.280 ;
        RECT 1126.730 0.010 1131.410 4.280 ;
        RECT 1132.250 0.010 1136.930 4.280 ;
        RECT 1137.770 0.010 1142.450 4.280 ;
        RECT 1143.290 0.010 1147.510 4.280 ;
        RECT 1148.350 0.010 1153.030 4.280 ;
        RECT 1153.870 0.010 1158.550 4.280 ;
        RECT 1159.390 0.010 1164.070 4.280 ;
        RECT 1164.910 0.010 1169.130 4.280 ;
        RECT 1169.970 0.010 1174.650 4.280 ;
        RECT 1175.490 0.010 1180.170 4.280 ;
        RECT 1181.010 0.010 1185.690 4.280 ;
        RECT 1186.530 0.010 1190.750 4.280 ;
        RECT 1191.590 0.010 1196.270 4.280 ;
        RECT 1197.110 0.010 1201.790 4.280 ;
        RECT 1202.630 0.010 1207.310 4.280 ;
        RECT 1208.150 0.010 1212.370 4.280 ;
        RECT 1213.210 0.010 1217.890 4.280 ;
        RECT 1218.730 0.010 1223.410 4.280 ;
        RECT 1224.250 0.010 1228.930 4.280 ;
        RECT 1229.770 0.010 1233.990 4.280 ;
        RECT 1234.830 0.010 1239.510 4.280 ;
        RECT 1240.350 0.010 1245.030 4.280 ;
        RECT 1245.870 0.010 1250.550 4.280 ;
        RECT 1251.390 0.010 1255.610 4.280 ;
        RECT 1256.450 0.010 1261.130 4.280 ;
        RECT 1261.970 0.010 1266.650 4.280 ;
        RECT 1267.490 0.010 1272.170 4.280 ;
        RECT 1273.010 0.010 1277.230 4.280 ;
        RECT 1278.070 0.010 1282.750 4.280 ;
        RECT 1283.590 0.010 1288.270 4.280 ;
        RECT 1289.110 0.010 1293.790 4.280 ;
        RECT 1294.630 0.010 1298.850 4.280 ;
        RECT 1299.690 0.010 1304.370 4.280 ;
        RECT 1305.210 0.010 1309.890 4.280 ;
        RECT 1310.730 0.010 1315.410 4.280 ;
        RECT 1316.250 0.010 1320.470 4.280 ;
        RECT 1321.310 0.010 1325.990 4.280 ;
        RECT 1326.830 0.010 1331.510 4.280 ;
        RECT 1332.350 0.010 1337.030 4.280 ;
        RECT 1337.870 0.010 1342.090 4.280 ;
        RECT 1342.930 0.010 1347.610 4.280 ;
        RECT 1348.450 0.010 1353.130 4.280 ;
        RECT 1353.970 0.010 1358.650 4.280 ;
        RECT 1359.490 0.010 1363.710 4.280 ;
        RECT 1364.550 0.010 1369.230 4.280 ;
        RECT 1370.070 0.010 1374.750 4.280 ;
        RECT 1375.590 0.010 1380.270 4.280 ;
        RECT 1381.110 0.010 1385.330 4.280 ;
        RECT 1386.170 0.010 1390.850 4.280 ;
        RECT 1391.690 0.010 1396.370 4.280 ;
      LAYER met3 ;
        RECT 4.400 1498.360 1377.175 1499.225 ;
        RECT 0.270 1497.720 1377.175 1498.360 ;
        RECT 4.400 1494.960 1377.175 1497.720 ;
        RECT 0.270 1494.320 1377.175 1494.960 ;
        RECT 4.400 1492.920 1377.175 1494.320 ;
        RECT 0.270 1492.280 1377.175 1492.920 ;
        RECT 4.400 1489.520 1377.175 1492.280 ;
        RECT 0.270 1488.880 1377.175 1489.520 ;
        RECT 4.400 1487.480 1377.175 1488.880 ;
        RECT 0.270 1486.840 1377.175 1487.480 ;
        RECT 4.400 1484.080 1377.175 1486.840 ;
        RECT 0.270 1483.440 1377.175 1484.080 ;
        RECT 4.400 1480.680 1377.175 1483.440 ;
        RECT 0.270 1480.040 1377.175 1480.680 ;
        RECT 4.400 1478.640 1377.175 1480.040 ;
        RECT 0.270 1478.000 1377.175 1478.640 ;
        RECT 4.400 1475.240 1377.175 1478.000 ;
        RECT 0.270 1474.600 1377.175 1475.240 ;
        RECT 4.400 1473.200 1377.175 1474.600 ;
        RECT 0.270 1472.560 1377.175 1473.200 ;
        RECT 4.400 1469.800 1377.175 1472.560 ;
        RECT 0.270 1469.160 1377.175 1469.800 ;
        RECT 4.400 1466.400 1377.175 1469.160 ;
        RECT 0.270 1465.760 1377.175 1466.400 ;
        RECT 4.400 1464.360 1377.175 1465.760 ;
        RECT 0.270 1463.720 1377.175 1464.360 ;
        RECT 4.400 1460.960 1377.175 1463.720 ;
        RECT 0.270 1460.320 1377.175 1460.960 ;
        RECT 4.400 1458.920 1377.175 1460.320 ;
        RECT 0.270 1458.280 1377.175 1458.920 ;
        RECT 4.400 1455.520 1377.175 1458.280 ;
        RECT 0.270 1454.880 1377.175 1455.520 ;
        RECT 4.400 1452.120 1377.175 1454.880 ;
        RECT 0.270 1451.480 1377.175 1452.120 ;
        RECT 4.400 1450.080 1377.175 1451.480 ;
        RECT 0.270 1449.440 1377.175 1450.080 ;
        RECT 4.400 1446.680 1377.175 1449.440 ;
        RECT 0.270 1446.040 1377.175 1446.680 ;
        RECT 4.400 1444.640 1377.175 1446.040 ;
        RECT 0.270 1444.000 1377.175 1444.640 ;
        RECT 4.400 1441.240 1377.175 1444.000 ;
        RECT 0.270 1440.600 1377.175 1441.240 ;
        RECT 4.400 1437.840 1377.175 1440.600 ;
        RECT 0.270 1437.200 1377.175 1437.840 ;
        RECT 4.400 1435.800 1377.175 1437.200 ;
        RECT 0.270 1435.160 1377.175 1435.800 ;
        RECT 4.400 1432.400 1377.175 1435.160 ;
        RECT 0.270 1431.760 1377.175 1432.400 ;
        RECT 4.400 1430.360 1377.175 1431.760 ;
        RECT 0.270 1429.720 1377.175 1430.360 ;
        RECT 4.400 1426.960 1377.175 1429.720 ;
        RECT 0.270 1426.320 1377.175 1426.960 ;
        RECT 4.400 1423.560 1377.175 1426.320 ;
        RECT 0.270 1422.920 1377.175 1423.560 ;
        RECT 4.400 1421.520 1377.175 1422.920 ;
        RECT 0.270 1420.880 1377.175 1421.520 ;
        RECT 4.400 1418.120 1377.175 1420.880 ;
        RECT 0.270 1417.480 1377.175 1418.120 ;
        RECT 4.400 1416.080 1377.175 1417.480 ;
        RECT 0.270 1415.440 1377.175 1416.080 ;
        RECT 4.400 1412.680 1377.175 1415.440 ;
        RECT 0.270 1412.040 1377.175 1412.680 ;
        RECT 4.400 1409.280 1377.175 1412.040 ;
        RECT 0.270 1408.640 1377.175 1409.280 ;
        RECT 4.400 1407.240 1377.175 1408.640 ;
        RECT 0.270 1406.600 1377.175 1407.240 ;
        RECT 4.400 1403.840 1377.175 1406.600 ;
        RECT 0.270 1403.200 1377.175 1403.840 ;
        RECT 4.400 1401.800 1377.175 1403.200 ;
        RECT 0.270 1401.160 1377.175 1401.800 ;
        RECT 4.400 1398.400 1377.175 1401.160 ;
        RECT 0.270 1397.760 1377.175 1398.400 ;
        RECT 4.400 1395.000 1377.175 1397.760 ;
        RECT 0.270 1394.360 1377.175 1395.000 ;
        RECT 4.400 1392.960 1377.175 1394.360 ;
        RECT 0.270 1392.320 1377.175 1392.960 ;
        RECT 4.400 1389.560 1377.175 1392.320 ;
        RECT 0.270 1388.920 1377.175 1389.560 ;
        RECT 4.400 1387.520 1377.175 1388.920 ;
        RECT 0.270 1386.880 1377.175 1387.520 ;
        RECT 4.400 1384.120 1377.175 1386.880 ;
        RECT 0.270 1383.480 1377.175 1384.120 ;
        RECT 4.400 1380.720 1377.175 1383.480 ;
        RECT 0.270 1380.080 1377.175 1380.720 ;
        RECT 4.400 1378.680 1377.175 1380.080 ;
        RECT 0.270 1378.040 1377.175 1378.680 ;
        RECT 4.400 1375.280 1377.175 1378.040 ;
        RECT 0.270 1374.640 1377.175 1375.280 ;
        RECT 4.400 1373.240 1377.175 1374.640 ;
        RECT 0.270 1372.600 1377.175 1373.240 ;
        RECT 4.400 1369.840 1377.175 1372.600 ;
        RECT 0.270 1369.200 1377.175 1369.840 ;
        RECT 4.400 1366.440 1377.175 1369.200 ;
        RECT 0.270 1365.800 1377.175 1366.440 ;
        RECT 4.400 1364.400 1377.175 1365.800 ;
        RECT 0.270 1363.760 1377.175 1364.400 ;
        RECT 4.400 1361.000 1377.175 1363.760 ;
        RECT 0.270 1360.360 1377.175 1361.000 ;
        RECT 4.400 1358.960 1377.175 1360.360 ;
        RECT 0.270 1358.320 1377.175 1358.960 ;
        RECT 4.400 1355.560 1377.175 1358.320 ;
        RECT 0.270 1354.920 1377.175 1355.560 ;
        RECT 4.400 1352.160 1377.175 1354.920 ;
        RECT 0.270 1351.520 1377.175 1352.160 ;
        RECT 4.400 1350.120 1377.175 1351.520 ;
        RECT 0.270 1349.480 1377.175 1350.120 ;
        RECT 4.400 1346.720 1377.175 1349.480 ;
        RECT 0.270 1346.080 1377.175 1346.720 ;
        RECT 4.400 1344.680 1377.175 1346.080 ;
        RECT 0.270 1344.040 1377.175 1344.680 ;
        RECT 4.400 1341.280 1377.175 1344.040 ;
        RECT 0.270 1340.640 1377.175 1341.280 ;
        RECT 4.400 1337.880 1377.175 1340.640 ;
        RECT 0.270 1337.240 1377.175 1337.880 ;
        RECT 4.400 1335.840 1377.175 1337.240 ;
        RECT 0.270 1335.200 1377.175 1335.840 ;
        RECT 4.400 1332.440 1377.175 1335.200 ;
        RECT 0.270 1331.800 1377.175 1332.440 ;
        RECT 4.400 1330.400 1377.175 1331.800 ;
        RECT 0.270 1329.760 1377.175 1330.400 ;
        RECT 4.400 1327.000 1377.175 1329.760 ;
        RECT 0.270 1326.360 1377.175 1327.000 ;
        RECT 4.400 1323.600 1377.175 1326.360 ;
        RECT 0.270 1322.960 1377.175 1323.600 ;
        RECT 4.400 1321.560 1377.175 1322.960 ;
        RECT 0.270 1320.920 1377.175 1321.560 ;
        RECT 4.400 1318.160 1377.175 1320.920 ;
        RECT 0.270 1317.520 1377.175 1318.160 ;
        RECT 4.400 1316.120 1377.175 1317.520 ;
        RECT 0.270 1315.480 1377.175 1316.120 ;
        RECT 4.400 1312.720 1377.175 1315.480 ;
        RECT 0.270 1312.080 1377.175 1312.720 ;
        RECT 4.400 1310.680 1377.175 1312.080 ;
        RECT 0.270 1310.040 1377.175 1310.680 ;
        RECT 4.400 1307.280 1377.175 1310.040 ;
        RECT 0.270 1306.640 1377.175 1307.280 ;
        RECT 4.400 1303.880 1377.175 1306.640 ;
        RECT 0.270 1303.240 1377.175 1303.880 ;
        RECT 4.400 1301.840 1377.175 1303.240 ;
        RECT 0.270 1301.200 1377.175 1301.840 ;
        RECT 4.400 1298.440 1377.175 1301.200 ;
        RECT 0.270 1297.800 1377.175 1298.440 ;
        RECT 4.400 1296.400 1377.175 1297.800 ;
        RECT 0.270 1295.760 1377.175 1296.400 ;
        RECT 4.400 1293.000 1377.175 1295.760 ;
        RECT 0.270 1292.360 1377.175 1293.000 ;
        RECT 4.400 1289.600 1377.175 1292.360 ;
        RECT 0.270 1288.960 1377.175 1289.600 ;
        RECT 4.400 1287.560 1377.175 1288.960 ;
        RECT 0.270 1286.920 1377.175 1287.560 ;
        RECT 4.400 1284.160 1377.175 1286.920 ;
        RECT 0.270 1283.520 1377.175 1284.160 ;
        RECT 4.400 1282.120 1377.175 1283.520 ;
        RECT 0.270 1281.480 1377.175 1282.120 ;
        RECT 4.400 1278.720 1377.175 1281.480 ;
        RECT 0.270 1278.080 1377.175 1278.720 ;
        RECT 4.400 1275.320 1377.175 1278.080 ;
        RECT 0.270 1274.680 1377.175 1275.320 ;
        RECT 4.400 1273.280 1377.175 1274.680 ;
        RECT 0.270 1272.640 1377.175 1273.280 ;
        RECT 4.400 1269.880 1377.175 1272.640 ;
        RECT 0.270 1269.240 1377.175 1269.880 ;
        RECT 4.400 1267.840 1377.175 1269.240 ;
        RECT 0.270 1267.200 1377.175 1267.840 ;
        RECT 4.400 1264.440 1377.175 1267.200 ;
        RECT 0.270 1263.800 1377.175 1264.440 ;
        RECT 4.400 1261.040 1377.175 1263.800 ;
        RECT 0.270 1260.400 1377.175 1261.040 ;
        RECT 4.400 1259.000 1377.175 1260.400 ;
        RECT 0.270 1258.360 1377.175 1259.000 ;
        RECT 4.400 1255.600 1377.175 1258.360 ;
        RECT 0.270 1254.960 1377.175 1255.600 ;
        RECT 4.400 1253.560 1377.175 1254.960 ;
        RECT 0.270 1252.920 1377.175 1253.560 ;
        RECT 4.400 1250.160 1377.175 1252.920 ;
        RECT 0.270 1249.520 1377.175 1250.160 ;
        RECT 4.400 1246.760 1377.175 1249.520 ;
        RECT 0.270 1246.120 1377.175 1246.760 ;
        RECT 4.400 1244.720 1377.175 1246.120 ;
        RECT 0.270 1244.080 1377.175 1244.720 ;
        RECT 4.400 1241.320 1377.175 1244.080 ;
        RECT 0.270 1240.680 1377.175 1241.320 ;
        RECT 4.400 1239.280 1377.175 1240.680 ;
        RECT 0.270 1238.640 1377.175 1239.280 ;
        RECT 4.400 1235.880 1377.175 1238.640 ;
        RECT 0.270 1235.240 1377.175 1235.880 ;
        RECT 4.400 1232.480 1377.175 1235.240 ;
        RECT 0.270 1231.840 1377.175 1232.480 ;
        RECT 4.400 1230.440 1377.175 1231.840 ;
        RECT 0.270 1229.800 1377.175 1230.440 ;
        RECT 4.400 1227.040 1377.175 1229.800 ;
        RECT 0.270 1226.400 1377.175 1227.040 ;
        RECT 4.400 1225.000 1377.175 1226.400 ;
        RECT 0.270 1224.360 1377.175 1225.000 ;
        RECT 4.400 1221.600 1377.175 1224.360 ;
        RECT 0.270 1220.960 1377.175 1221.600 ;
        RECT 4.400 1218.200 1377.175 1220.960 ;
        RECT 0.270 1217.560 1377.175 1218.200 ;
        RECT 4.400 1216.160 1377.175 1217.560 ;
        RECT 0.270 1215.520 1377.175 1216.160 ;
        RECT 4.400 1212.760 1377.175 1215.520 ;
        RECT 0.270 1212.120 1377.175 1212.760 ;
        RECT 4.400 1210.720 1377.175 1212.120 ;
        RECT 0.270 1210.080 1377.175 1210.720 ;
        RECT 4.400 1207.320 1377.175 1210.080 ;
        RECT 0.270 1206.680 1377.175 1207.320 ;
        RECT 4.400 1203.920 1377.175 1206.680 ;
        RECT 0.270 1203.280 1377.175 1203.920 ;
        RECT 4.400 1201.880 1377.175 1203.280 ;
        RECT 0.270 1201.240 1377.175 1201.880 ;
        RECT 4.400 1198.480 1377.175 1201.240 ;
        RECT 0.270 1197.840 1377.175 1198.480 ;
        RECT 4.400 1196.440 1377.175 1197.840 ;
        RECT 0.270 1195.800 1377.175 1196.440 ;
        RECT 4.400 1193.040 1377.175 1195.800 ;
        RECT 0.270 1192.400 1377.175 1193.040 ;
        RECT 4.400 1189.640 1377.175 1192.400 ;
        RECT 0.270 1189.000 1377.175 1189.640 ;
        RECT 4.400 1187.600 1377.175 1189.000 ;
        RECT 0.270 1186.960 1377.175 1187.600 ;
        RECT 4.400 1184.200 1377.175 1186.960 ;
        RECT 0.270 1183.560 1377.175 1184.200 ;
        RECT 4.400 1182.160 1377.175 1183.560 ;
        RECT 0.270 1181.520 1377.175 1182.160 ;
        RECT 4.400 1178.760 1377.175 1181.520 ;
        RECT 0.270 1178.120 1377.175 1178.760 ;
        RECT 4.400 1175.360 1377.175 1178.120 ;
        RECT 0.270 1174.720 1377.175 1175.360 ;
        RECT 4.400 1173.320 1377.175 1174.720 ;
        RECT 0.270 1172.680 1377.175 1173.320 ;
        RECT 4.400 1169.920 1377.175 1172.680 ;
        RECT 0.270 1169.280 1377.175 1169.920 ;
        RECT 4.400 1167.880 1377.175 1169.280 ;
        RECT 0.270 1167.240 1377.175 1167.880 ;
        RECT 4.400 1164.480 1377.175 1167.240 ;
        RECT 0.270 1163.840 1377.175 1164.480 ;
        RECT 4.400 1161.080 1377.175 1163.840 ;
        RECT 0.270 1160.440 1377.175 1161.080 ;
        RECT 4.400 1159.040 1377.175 1160.440 ;
        RECT 0.270 1158.400 1377.175 1159.040 ;
        RECT 4.400 1155.640 1377.175 1158.400 ;
        RECT 0.270 1155.000 1377.175 1155.640 ;
        RECT 4.400 1153.600 1377.175 1155.000 ;
        RECT 0.270 1152.960 1377.175 1153.600 ;
        RECT 4.400 1150.200 1377.175 1152.960 ;
        RECT 0.270 1149.560 1377.175 1150.200 ;
        RECT 4.400 1146.800 1377.175 1149.560 ;
        RECT 0.270 1146.160 1377.175 1146.800 ;
        RECT 4.400 1144.760 1377.175 1146.160 ;
        RECT 0.270 1144.120 1377.175 1144.760 ;
        RECT 4.400 1141.360 1377.175 1144.120 ;
        RECT 0.270 1140.720 1377.175 1141.360 ;
        RECT 4.400 1139.320 1377.175 1140.720 ;
        RECT 0.270 1138.680 1377.175 1139.320 ;
        RECT 4.400 1135.920 1377.175 1138.680 ;
        RECT 0.270 1135.280 1377.175 1135.920 ;
        RECT 4.400 1132.520 1377.175 1135.280 ;
        RECT 0.270 1131.880 1377.175 1132.520 ;
        RECT 4.400 1130.480 1377.175 1131.880 ;
        RECT 0.270 1129.840 1377.175 1130.480 ;
        RECT 4.400 1127.080 1377.175 1129.840 ;
        RECT 0.270 1126.440 1377.175 1127.080 ;
        RECT 4.400 1125.040 1377.175 1126.440 ;
        RECT 0.270 1124.400 1377.175 1125.040 ;
        RECT 4.400 1121.640 1377.175 1124.400 ;
        RECT 0.270 1121.000 1377.175 1121.640 ;
        RECT 4.400 1119.600 1377.175 1121.000 ;
        RECT 0.270 1118.960 1377.175 1119.600 ;
        RECT 4.400 1116.200 1377.175 1118.960 ;
        RECT 0.270 1115.560 1377.175 1116.200 ;
        RECT 4.400 1112.800 1377.175 1115.560 ;
        RECT 0.270 1112.160 1377.175 1112.800 ;
        RECT 4.400 1110.760 1377.175 1112.160 ;
        RECT 0.270 1110.120 1377.175 1110.760 ;
        RECT 4.400 1107.360 1377.175 1110.120 ;
        RECT 0.270 1106.720 1377.175 1107.360 ;
        RECT 4.400 1105.320 1377.175 1106.720 ;
        RECT 0.270 1104.680 1377.175 1105.320 ;
        RECT 4.400 1101.920 1377.175 1104.680 ;
        RECT 0.270 1101.280 1377.175 1101.920 ;
        RECT 4.400 1098.520 1377.175 1101.280 ;
        RECT 0.270 1097.880 1377.175 1098.520 ;
        RECT 4.400 1096.480 1377.175 1097.880 ;
        RECT 0.270 1095.840 1377.175 1096.480 ;
        RECT 4.400 1093.080 1377.175 1095.840 ;
        RECT 0.270 1092.440 1377.175 1093.080 ;
        RECT 4.400 1091.040 1377.175 1092.440 ;
        RECT 0.270 1090.400 1377.175 1091.040 ;
        RECT 4.400 1087.640 1377.175 1090.400 ;
        RECT 0.270 1087.000 1377.175 1087.640 ;
        RECT 4.400 1084.240 1377.175 1087.000 ;
        RECT 0.270 1083.600 1377.175 1084.240 ;
        RECT 4.400 1082.200 1377.175 1083.600 ;
        RECT 0.270 1081.560 1377.175 1082.200 ;
        RECT 4.400 1078.800 1377.175 1081.560 ;
        RECT 0.270 1078.160 1377.175 1078.800 ;
        RECT 4.400 1076.760 1377.175 1078.160 ;
        RECT 0.270 1076.120 1377.175 1076.760 ;
        RECT 4.400 1073.360 1377.175 1076.120 ;
        RECT 0.270 1072.720 1377.175 1073.360 ;
        RECT 4.400 1069.960 1377.175 1072.720 ;
        RECT 0.270 1069.320 1377.175 1069.960 ;
        RECT 4.400 1067.920 1377.175 1069.320 ;
        RECT 0.270 1067.280 1377.175 1067.920 ;
        RECT 4.400 1064.520 1377.175 1067.280 ;
        RECT 0.270 1063.880 1377.175 1064.520 ;
        RECT 4.400 1062.480 1377.175 1063.880 ;
        RECT 0.270 1061.840 1377.175 1062.480 ;
        RECT 4.400 1059.080 1377.175 1061.840 ;
        RECT 0.270 1058.440 1377.175 1059.080 ;
        RECT 4.400 1055.680 1377.175 1058.440 ;
        RECT 0.270 1055.040 1377.175 1055.680 ;
        RECT 4.400 1053.640 1377.175 1055.040 ;
        RECT 0.270 1053.000 1377.175 1053.640 ;
        RECT 4.400 1050.240 1377.175 1053.000 ;
        RECT 0.270 1049.600 1377.175 1050.240 ;
        RECT 4.400 1048.200 1377.175 1049.600 ;
        RECT 0.270 1047.560 1377.175 1048.200 ;
        RECT 4.400 1044.800 1377.175 1047.560 ;
        RECT 0.270 1044.160 1377.175 1044.800 ;
        RECT 4.400 1041.400 1377.175 1044.160 ;
        RECT 0.270 1040.760 1377.175 1041.400 ;
        RECT 4.400 1039.360 1377.175 1040.760 ;
        RECT 0.270 1038.720 1377.175 1039.360 ;
        RECT 4.400 1035.960 1377.175 1038.720 ;
        RECT 0.270 1035.320 1377.175 1035.960 ;
        RECT 4.400 1033.920 1377.175 1035.320 ;
        RECT 0.270 1033.280 1377.175 1033.920 ;
        RECT 4.400 1030.520 1377.175 1033.280 ;
        RECT 0.270 1029.880 1377.175 1030.520 ;
        RECT 4.400 1027.120 1377.175 1029.880 ;
        RECT 0.270 1026.480 1377.175 1027.120 ;
        RECT 4.400 1025.080 1377.175 1026.480 ;
        RECT 0.270 1024.440 1377.175 1025.080 ;
        RECT 4.400 1021.680 1377.175 1024.440 ;
        RECT 0.270 1021.040 1377.175 1021.680 ;
        RECT 4.400 1019.640 1377.175 1021.040 ;
        RECT 0.270 1019.000 1377.175 1019.640 ;
        RECT 4.400 1016.240 1377.175 1019.000 ;
        RECT 0.270 1015.600 1377.175 1016.240 ;
        RECT 4.400 1012.840 1377.175 1015.600 ;
        RECT 0.270 1012.200 1377.175 1012.840 ;
        RECT 4.400 1010.800 1377.175 1012.200 ;
        RECT 0.270 1010.160 1377.175 1010.800 ;
        RECT 4.400 1007.400 1377.175 1010.160 ;
        RECT 0.270 1006.760 1377.175 1007.400 ;
        RECT 4.400 1005.360 1377.175 1006.760 ;
        RECT 0.270 1004.720 1377.175 1005.360 ;
        RECT 4.400 1001.960 1377.175 1004.720 ;
        RECT 0.270 1001.320 1377.175 1001.960 ;
        RECT 4.400 998.560 1377.175 1001.320 ;
        RECT 0.270 997.920 1377.175 998.560 ;
        RECT 4.400 996.520 1377.175 997.920 ;
        RECT 0.270 995.880 1377.175 996.520 ;
        RECT 4.400 993.120 1377.175 995.880 ;
        RECT 0.270 992.480 1377.175 993.120 ;
        RECT 4.400 991.080 1377.175 992.480 ;
        RECT 0.270 990.440 1377.175 991.080 ;
        RECT 4.400 987.680 1377.175 990.440 ;
        RECT 0.270 987.040 1377.175 987.680 ;
        RECT 4.400 984.280 1377.175 987.040 ;
        RECT 0.270 983.640 1377.175 984.280 ;
        RECT 4.400 982.240 1377.175 983.640 ;
        RECT 0.270 981.600 1377.175 982.240 ;
        RECT 4.400 978.840 1377.175 981.600 ;
        RECT 0.270 978.200 1377.175 978.840 ;
        RECT 4.400 976.800 1377.175 978.200 ;
        RECT 0.270 976.160 1377.175 976.800 ;
        RECT 4.400 973.400 1377.175 976.160 ;
        RECT 0.270 972.760 1377.175 973.400 ;
        RECT 4.400 970.000 1377.175 972.760 ;
        RECT 0.270 969.360 1377.175 970.000 ;
        RECT 4.400 967.960 1377.175 969.360 ;
        RECT 0.270 967.320 1377.175 967.960 ;
        RECT 4.400 964.560 1377.175 967.320 ;
        RECT 0.270 963.920 1377.175 964.560 ;
        RECT 4.400 962.520 1377.175 963.920 ;
        RECT 0.270 961.880 1377.175 962.520 ;
        RECT 4.400 959.120 1377.175 961.880 ;
        RECT 0.270 958.480 1377.175 959.120 ;
        RECT 4.400 955.720 1377.175 958.480 ;
        RECT 0.270 955.080 1377.175 955.720 ;
        RECT 4.400 953.680 1377.175 955.080 ;
        RECT 0.270 953.040 1377.175 953.680 ;
        RECT 4.400 950.280 1377.175 953.040 ;
        RECT 0.270 949.640 1377.175 950.280 ;
        RECT 4.400 948.240 1377.175 949.640 ;
        RECT 0.270 947.600 1377.175 948.240 ;
        RECT 4.400 944.840 1377.175 947.600 ;
        RECT 0.270 944.200 1377.175 944.840 ;
        RECT 4.400 941.440 1377.175 944.200 ;
        RECT 0.270 940.800 1377.175 941.440 ;
        RECT 4.400 939.400 1377.175 940.800 ;
        RECT 0.270 938.760 1377.175 939.400 ;
        RECT 4.400 936.000 1377.175 938.760 ;
        RECT 0.270 935.360 1377.175 936.000 ;
        RECT 4.400 933.960 1377.175 935.360 ;
        RECT 0.270 933.320 1377.175 933.960 ;
        RECT 4.400 930.560 1377.175 933.320 ;
        RECT 0.270 929.920 1377.175 930.560 ;
        RECT 4.400 928.520 1377.175 929.920 ;
        RECT 0.270 927.880 1377.175 928.520 ;
        RECT 4.400 925.120 1377.175 927.880 ;
        RECT 0.270 924.480 1377.175 925.120 ;
        RECT 4.400 921.720 1377.175 924.480 ;
        RECT 0.270 921.080 1377.175 921.720 ;
        RECT 4.400 919.680 1377.175 921.080 ;
        RECT 0.270 919.040 1377.175 919.680 ;
        RECT 4.400 916.280 1377.175 919.040 ;
        RECT 0.270 915.640 1377.175 916.280 ;
        RECT 4.400 914.240 1377.175 915.640 ;
        RECT 0.270 913.600 1377.175 914.240 ;
        RECT 4.400 910.840 1377.175 913.600 ;
        RECT 0.270 910.200 1377.175 910.840 ;
        RECT 4.400 907.440 1377.175 910.200 ;
        RECT 0.270 906.800 1377.175 907.440 ;
        RECT 4.400 905.400 1377.175 906.800 ;
        RECT 0.270 904.760 1377.175 905.400 ;
        RECT 4.400 902.000 1377.175 904.760 ;
        RECT 0.270 901.360 1377.175 902.000 ;
        RECT 4.400 899.960 1377.175 901.360 ;
        RECT 0.270 899.320 1377.175 899.960 ;
        RECT 4.400 896.560 1377.175 899.320 ;
        RECT 0.270 895.920 1377.175 896.560 ;
        RECT 4.400 893.160 1377.175 895.920 ;
        RECT 0.270 892.520 1377.175 893.160 ;
        RECT 4.400 891.120 1377.175 892.520 ;
        RECT 0.270 890.480 1377.175 891.120 ;
        RECT 4.400 887.720 1377.175 890.480 ;
        RECT 0.270 887.080 1377.175 887.720 ;
        RECT 4.400 885.680 1377.175 887.080 ;
        RECT 0.270 885.040 1377.175 885.680 ;
        RECT 4.400 882.280 1377.175 885.040 ;
        RECT 0.270 881.640 1377.175 882.280 ;
        RECT 4.400 878.880 1377.175 881.640 ;
        RECT 0.270 878.240 1377.175 878.880 ;
        RECT 4.400 876.840 1377.175 878.240 ;
        RECT 0.270 876.200 1377.175 876.840 ;
        RECT 4.400 873.440 1377.175 876.200 ;
        RECT 0.270 872.800 1377.175 873.440 ;
        RECT 4.400 871.400 1377.175 872.800 ;
        RECT 0.270 870.760 1377.175 871.400 ;
        RECT 4.400 868.000 1377.175 870.760 ;
        RECT 0.270 867.360 1377.175 868.000 ;
        RECT 4.400 864.600 1377.175 867.360 ;
        RECT 0.270 863.960 1377.175 864.600 ;
        RECT 4.400 862.560 1377.175 863.960 ;
        RECT 0.270 861.920 1377.175 862.560 ;
        RECT 4.400 859.160 1377.175 861.920 ;
        RECT 0.270 858.520 1377.175 859.160 ;
        RECT 4.400 857.120 1377.175 858.520 ;
        RECT 0.270 856.480 1377.175 857.120 ;
        RECT 4.400 853.720 1377.175 856.480 ;
        RECT 0.270 853.080 1377.175 853.720 ;
        RECT 4.400 850.320 1377.175 853.080 ;
        RECT 0.270 849.680 1377.175 850.320 ;
        RECT 4.400 848.280 1377.175 849.680 ;
        RECT 0.270 847.640 1377.175 848.280 ;
        RECT 4.400 844.880 1377.175 847.640 ;
        RECT 0.270 844.240 1377.175 844.880 ;
        RECT 4.400 842.840 1377.175 844.240 ;
        RECT 0.270 842.200 1377.175 842.840 ;
        RECT 4.400 839.440 1377.175 842.200 ;
        RECT 0.270 838.800 1377.175 839.440 ;
        RECT 4.400 836.040 1377.175 838.800 ;
        RECT 0.270 835.400 1377.175 836.040 ;
        RECT 4.400 834.000 1377.175 835.400 ;
        RECT 0.270 833.360 1377.175 834.000 ;
        RECT 4.400 830.600 1377.175 833.360 ;
        RECT 0.270 829.960 1377.175 830.600 ;
        RECT 4.400 828.560 1377.175 829.960 ;
        RECT 0.270 827.920 1377.175 828.560 ;
        RECT 4.400 825.160 1377.175 827.920 ;
        RECT 0.270 824.520 1377.175 825.160 ;
        RECT 4.400 821.760 1377.175 824.520 ;
        RECT 0.270 821.120 1377.175 821.760 ;
        RECT 4.400 819.720 1377.175 821.120 ;
        RECT 0.270 819.080 1377.175 819.720 ;
        RECT 4.400 816.320 1377.175 819.080 ;
        RECT 0.270 815.680 1377.175 816.320 ;
        RECT 4.400 814.280 1377.175 815.680 ;
        RECT 0.270 813.640 1377.175 814.280 ;
        RECT 4.400 810.880 1377.175 813.640 ;
        RECT 0.270 810.240 1377.175 810.880 ;
        RECT 4.400 807.480 1377.175 810.240 ;
        RECT 0.270 806.840 1377.175 807.480 ;
        RECT 4.400 805.440 1377.175 806.840 ;
        RECT 0.270 804.800 1377.175 805.440 ;
        RECT 4.400 802.040 1377.175 804.800 ;
        RECT 0.270 801.400 1377.175 802.040 ;
        RECT 4.400 800.000 1377.175 801.400 ;
        RECT 0.270 799.360 1377.175 800.000 ;
        RECT 4.400 796.600 1377.175 799.360 ;
        RECT 0.270 795.960 1377.175 796.600 ;
        RECT 4.400 793.200 1377.175 795.960 ;
        RECT 0.270 792.560 1377.175 793.200 ;
        RECT 4.400 791.160 1377.175 792.560 ;
        RECT 0.270 790.520 1377.175 791.160 ;
        RECT 4.400 787.760 1377.175 790.520 ;
        RECT 0.270 787.120 1377.175 787.760 ;
        RECT 4.400 785.720 1377.175 787.120 ;
        RECT 0.270 785.080 1377.175 785.720 ;
        RECT 4.400 782.320 1377.175 785.080 ;
        RECT 0.270 781.680 1377.175 782.320 ;
        RECT 4.400 778.920 1377.175 781.680 ;
        RECT 0.270 778.280 1377.175 778.920 ;
        RECT 4.400 776.880 1377.175 778.280 ;
        RECT 0.270 776.240 1377.175 776.880 ;
        RECT 4.400 773.480 1377.175 776.240 ;
        RECT 0.270 772.840 1377.175 773.480 ;
        RECT 4.400 771.440 1377.175 772.840 ;
        RECT 0.270 770.800 1377.175 771.440 ;
        RECT 4.400 768.040 1377.175 770.800 ;
        RECT 0.270 767.400 1377.175 768.040 ;
        RECT 4.400 764.640 1377.175 767.400 ;
        RECT 0.270 764.000 1377.175 764.640 ;
        RECT 4.400 762.600 1377.175 764.000 ;
        RECT 0.270 761.960 1377.175 762.600 ;
        RECT 4.400 759.200 1377.175 761.960 ;
        RECT 0.270 758.560 1377.175 759.200 ;
        RECT 4.400 757.160 1377.175 758.560 ;
        RECT 0.270 756.520 1377.175 757.160 ;
        RECT 4.400 753.760 1377.175 756.520 ;
        RECT 0.270 753.120 1377.175 753.760 ;
        RECT 4.400 750.360 1377.175 753.120 ;
        RECT 0.270 749.720 1377.175 750.360 ;
        RECT 4.400 748.320 1377.175 749.720 ;
        RECT 0.270 747.680 1377.175 748.320 ;
        RECT 4.400 744.920 1377.175 747.680 ;
        RECT 0.270 744.280 1377.175 744.920 ;
        RECT 4.400 742.880 1377.175 744.280 ;
        RECT 0.270 742.240 1377.175 742.880 ;
        RECT 4.400 739.480 1377.175 742.240 ;
        RECT 0.270 738.840 1377.175 739.480 ;
        RECT 4.400 737.440 1377.175 738.840 ;
        RECT 0.270 736.800 1377.175 737.440 ;
        RECT 4.400 734.040 1377.175 736.800 ;
        RECT 0.270 733.400 1377.175 734.040 ;
        RECT 4.400 730.640 1377.175 733.400 ;
        RECT 0.270 730.000 1377.175 730.640 ;
        RECT 4.400 728.600 1377.175 730.000 ;
        RECT 0.270 727.960 1377.175 728.600 ;
        RECT 4.400 725.200 1377.175 727.960 ;
        RECT 0.270 724.560 1377.175 725.200 ;
        RECT 4.400 723.160 1377.175 724.560 ;
        RECT 0.270 722.520 1377.175 723.160 ;
        RECT 4.400 719.760 1377.175 722.520 ;
        RECT 0.270 719.120 1377.175 719.760 ;
        RECT 4.400 716.360 1377.175 719.120 ;
        RECT 0.270 715.720 1377.175 716.360 ;
        RECT 4.400 714.320 1377.175 715.720 ;
        RECT 0.270 713.680 1377.175 714.320 ;
        RECT 4.400 710.920 1377.175 713.680 ;
        RECT 0.270 710.280 1377.175 710.920 ;
        RECT 4.400 708.880 1377.175 710.280 ;
        RECT 0.270 708.240 1377.175 708.880 ;
        RECT 4.400 705.480 1377.175 708.240 ;
        RECT 0.270 704.840 1377.175 705.480 ;
        RECT 4.400 702.080 1377.175 704.840 ;
        RECT 0.270 701.440 1377.175 702.080 ;
        RECT 4.400 700.040 1377.175 701.440 ;
        RECT 0.270 699.400 1377.175 700.040 ;
        RECT 4.400 696.640 1377.175 699.400 ;
        RECT 0.270 696.000 1377.175 696.640 ;
        RECT 4.400 694.600 1377.175 696.000 ;
        RECT 0.270 693.960 1377.175 694.600 ;
        RECT 4.400 691.200 1377.175 693.960 ;
        RECT 0.270 690.560 1377.175 691.200 ;
        RECT 4.400 687.800 1377.175 690.560 ;
        RECT 0.270 687.160 1377.175 687.800 ;
        RECT 4.400 685.760 1377.175 687.160 ;
        RECT 0.270 685.120 1377.175 685.760 ;
        RECT 4.400 682.360 1377.175 685.120 ;
        RECT 0.270 681.720 1377.175 682.360 ;
        RECT 4.400 680.320 1377.175 681.720 ;
        RECT 0.270 679.680 1377.175 680.320 ;
        RECT 4.400 676.920 1377.175 679.680 ;
        RECT 0.270 676.280 1377.175 676.920 ;
        RECT 4.400 673.520 1377.175 676.280 ;
        RECT 0.270 672.880 1377.175 673.520 ;
        RECT 4.400 671.480 1377.175 672.880 ;
        RECT 0.270 670.840 1377.175 671.480 ;
        RECT 4.400 668.080 1377.175 670.840 ;
        RECT 0.270 667.440 1377.175 668.080 ;
        RECT 4.400 666.040 1377.175 667.440 ;
        RECT 0.270 665.400 1377.175 666.040 ;
        RECT 4.400 662.640 1377.175 665.400 ;
        RECT 0.270 662.000 1377.175 662.640 ;
        RECT 4.400 659.240 1377.175 662.000 ;
        RECT 0.270 658.600 1377.175 659.240 ;
        RECT 4.400 657.200 1377.175 658.600 ;
        RECT 0.270 656.560 1377.175 657.200 ;
        RECT 4.400 653.800 1377.175 656.560 ;
        RECT 0.270 653.160 1377.175 653.800 ;
        RECT 4.400 651.760 1377.175 653.160 ;
        RECT 0.270 651.120 1377.175 651.760 ;
        RECT 4.400 648.360 1377.175 651.120 ;
        RECT 0.270 647.720 1377.175 648.360 ;
        RECT 4.400 644.960 1377.175 647.720 ;
        RECT 0.270 644.320 1377.175 644.960 ;
        RECT 4.400 642.920 1377.175 644.320 ;
        RECT 0.270 642.280 1377.175 642.920 ;
        RECT 4.400 639.520 1377.175 642.280 ;
        RECT 0.270 638.880 1377.175 639.520 ;
        RECT 4.400 637.480 1377.175 638.880 ;
        RECT 0.270 636.840 1377.175 637.480 ;
        RECT 4.400 634.080 1377.175 636.840 ;
        RECT 0.270 633.440 1377.175 634.080 ;
        RECT 4.400 630.680 1377.175 633.440 ;
        RECT 0.270 630.040 1377.175 630.680 ;
        RECT 4.400 628.640 1377.175 630.040 ;
        RECT 0.270 628.000 1377.175 628.640 ;
        RECT 4.400 625.240 1377.175 628.000 ;
        RECT 0.270 624.600 1377.175 625.240 ;
        RECT 4.400 623.200 1377.175 624.600 ;
        RECT 0.270 622.560 1377.175 623.200 ;
        RECT 4.400 619.800 1377.175 622.560 ;
        RECT 0.270 619.160 1377.175 619.800 ;
        RECT 4.400 616.400 1377.175 619.160 ;
        RECT 0.270 615.760 1377.175 616.400 ;
        RECT 4.400 614.360 1377.175 615.760 ;
        RECT 0.270 613.720 1377.175 614.360 ;
        RECT 4.400 610.960 1377.175 613.720 ;
        RECT 0.270 610.320 1377.175 610.960 ;
        RECT 4.400 608.920 1377.175 610.320 ;
        RECT 0.270 608.280 1377.175 608.920 ;
        RECT 4.400 605.520 1377.175 608.280 ;
        RECT 0.270 604.880 1377.175 605.520 ;
        RECT 4.400 602.120 1377.175 604.880 ;
        RECT 0.270 601.480 1377.175 602.120 ;
        RECT 4.400 600.080 1377.175 601.480 ;
        RECT 0.270 599.440 1377.175 600.080 ;
        RECT 4.400 596.680 1377.175 599.440 ;
        RECT 0.270 596.040 1377.175 596.680 ;
        RECT 4.400 594.640 1377.175 596.040 ;
        RECT 0.270 594.000 1377.175 594.640 ;
        RECT 4.400 591.240 1377.175 594.000 ;
        RECT 0.270 590.600 1377.175 591.240 ;
        RECT 4.400 587.840 1377.175 590.600 ;
        RECT 0.270 587.200 1377.175 587.840 ;
        RECT 4.400 585.800 1377.175 587.200 ;
        RECT 0.270 585.160 1377.175 585.800 ;
        RECT 4.400 582.400 1377.175 585.160 ;
        RECT 0.270 581.760 1377.175 582.400 ;
        RECT 4.400 580.360 1377.175 581.760 ;
        RECT 0.270 579.720 1377.175 580.360 ;
        RECT 4.400 576.960 1377.175 579.720 ;
        RECT 0.270 576.320 1377.175 576.960 ;
        RECT 4.400 573.560 1377.175 576.320 ;
        RECT 0.270 572.920 1377.175 573.560 ;
        RECT 4.400 571.520 1377.175 572.920 ;
        RECT 0.270 570.880 1377.175 571.520 ;
        RECT 4.400 568.120 1377.175 570.880 ;
        RECT 0.270 567.480 1377.175 568.120 ;
        RECT 4.400 566.080 1377.175 567.480 ;
        RECT 0.270 565.440 1377.175 566.080 ;
        RECT 4.400 562.680 1377.175 565.440 ;
        RECT 0.270 562.040 1377.175 562.680 ;
        RECT 4.400 560.640 1377.175 562.040 ;
        RECT 0.270 560.000 1377.175 560.640 ;
        RECT 4.400 557.240 1377.175 560.000 ;
        RECT 0.270 556.600 1377.175 557.240 ;
        RECT 4.400 553.840 1377.175 556.600 ;
        RECT 0.270 553.200 1377.175 553.840 ;
        RECT 4.400 551.800 1377.175 553.200 ;
        RECT 0.270 551.160 1377.175 551.800 ;
        RECT 4.400 548.400 1377.175 551.160 ;
        RECT 0.270 547.760 1377.175 548.400 ;
        RECT 4.400 546.360 1377.175 547.760 ;
        RECT 0.270 545.720 1377.175 546.360 ;
        RECT 4.400 542.960 1377.175 545.720 ;
        RECT 0.270 542.320 1377.175 542.960 ;
        RECT 4.400 539.560 1377.175 542.320 ;
        RECT 0.270 538.920 1377.175 539.560 ;
        RECT 4.400 537.520 1377.175 538.920 ;
        RECT 0.270 536.880 1377.175 537.520 ;
        RECT 4.400 534.120 1377.175 536.880 ;
        RECT 0.270 533.480 1377.175 534.120 ;
        RECT 4.400 532.080 1377.175 533.480 ;
        RECT 0.270 531.440 1377.175 532.080 ;
        RECT 4.400 528.680 1377.175 531.440 ;
        RECT 0.270 528.040 1377.175 528.680 ;
        RECT 4.400 525.280 1377.175 528.040 ;
        RECT 0.270 524.640 1377.175 525.280 ;
        RECT 4.400 523.240 1377.175 524.640 ;
        RECT 0.270 522.600 1377.175 523.240 ;
        RECT 4.400 519.840 1377.175 522.600 ;
        RECT 0.270 519.200 1377.175 519.840 ;
        RECT 4.400 517.800 1377.175 519.200 ;
        RECT 0.270 517.160 1377.175 517.800 ;
        RECT 4.400 514.400 1377.175 517.160 ;
        RECT 0.270 513.760 1377.175 514.400 ;
        RECT 4.400 511.000 1377.175 513.760 ;
        RECT 0.270 510.360 1377.175 511.000 ;
        RECT 4.400 508.960 1377.175 510.360 ;
        RECT 0.270 508.320 1377.175 508.960 ;
        RECT 4.400 505.560 1377.175 508.320 ;
        RECT 0.270 504.920 1377.175 505.560 ;
        RECT 4.400 503.520 1377.175 504.920 ;
        RECT 0.270 502.880 1377.175 503.520 ;
        RECT 4.400 500.120 1377.175 502.880 ;
        RECT 0.270 499.480 1377.175 500.120 ;
        RECT 4.400 496.720 1377.175 499.480 ;
        RECT 0.270 496.080 1377.175 496.720 ;
        RECT 4.400 494.680 1377.175 496.080 ;
        RECT 0.270 494.040 1377.175 494.680 ;
        RECT 4.400 491.280 1377.175 494.040 ;
        RECT 0.270 490.640 1377.175 491.280 ;
        RECT 4.400 489.240 1377.175 490.640 ;
        RECT 0.270 488.600 1377.175 489.240 ;
        RECT 4.400 485.840 1377.175 488.600 ;
        RECT 0.270 485.200 1377.175 485.840 ;
        RECT 4.400 482.440 1377.175 485.200 ;
        RECT 0.270 481.800 1377.175 482.440 ;
        RECT 4.400 480.400 1377.175 481.800 ;
        RECT 0.270 479.760 1377.175 480.400 ;
        RECT 4.400 477.000 1377.175 479.760 ;
        RECT 0.270 476.360 1377.175 477.000 ;
        RECT 4.400 474.960 1377.175 476.360 ;
        RECT 0.270 474.320 1377.175 474.960 ;
        RECT 4.400 471.560 1377.175 474.320 ;
        RECT 0.270 470.920 1377.175 471.560 ;
        RECT 4.400 468.160 1377.175 470.920 ;
        RECT 0.270 467.520 1377.175 468.160 ;
        RECT 4.400 466.120 1377.175 467.520 ;
        RECT 0.270 465.480 1377.175 466.120 ;
        RECT 4.400 462.720 1377.175 465.480 ;
        RECT 0.270 462.080 1377.175 462.720 ;
        RECT 4.400 460.680 1377.175 462.080 ;
        RECT 0.270 460.040 1377.175 460.680 ;
        RECT 4.400 457.280 1377.175 460.040 ;
        RECT 0.270 456.640 1377.175 457.280 ;
        RECT 4.400 453.880 1377.175 456.640 ;
        RECT 0.270 453.240 1377.175 453.880 ;
        RECT 4.400 451.840 1377.175 453.240 ;
        RECT 0.270 451.200 1377.175 451.840 ;
        RECT 4.400 448.440 1377.175 451.200 ;
        RECT 0.270 447.800 1377.175 448.440 ;
        RECT 4.400 446.400 1377.175 447.800 ;
        RECT 0.270 445.760 1377.175 446.400 ;
        RECT 4.400 443.000 1377.175 445.760 ;
        RECT 0.270 442.360 1377.175 443.000 ;
        RECT 4.400 439.600 1377.175 442.360 ;
        RECT 0.270 438.960 1377.175 439.600 ;
        RECT 4.400 437.560 1377.175 438.960 ;
        RECT 0.270 436.920 1377.175 437.560 ;
        RECT 4.400 434.160 1377.175 436.920 ;
        RECT 0.270 433.520 1377.175 434.160 ;
        RECT 4.400 432.120 1377.175 433.520 ;
        RECT 0.270 431.480 1377.175 432.120 ;
        RECT 4.400 428.720 1377.175 431.480 ;
        RECT 0.270 428.080 1377.175 428.720 ;
        RECT 4.400 425.320 1377.175 428.080 ;
        RECT 0.270 424.680 1377.175 425.320 ;
        RECT 4.400 423.280 1377.175 424.680 ;
        RECT 0.270 422.640 1377.175 423.280 ;
        RECT 4.400 419.880 1377.175 422.640 ;
        RECT 0.270 419.240 1377.175 419.880 ;
        RECT 4.400 417.840 1377.175 419.240 ;
        RECT 0.270 417.200 1377.175 417.840 ;
        RECT 4.400 414.440 1377.175 417.200 ;
        RECT 0.270 413.800 1377.175 414.440 ;
        RECT 4.400 411.040 1377.175 413.800 ;
        RECT 0.270 410.400 1377.175 411.040 ;
        RECT 4.400 409.000 1377.175 410.400 ;
        RECT 0.270 408.360 1377.175 409.000 ;
        RECT 4.400 405.600 1377.175 408.360 ;
        RECT 0.270 404.960 1377.175 405.600 ;
        RECT 4.400 403.560 1377.175 404.960 ;
        RECT 0.270 402.920 1377.175 403.560 ;
        RECT 4.400 400.160 1377.175 402.920 ;
        RECT 0.270 399.520 1377.175 400.160 ;
        RECT 4.400 396.760 1377.175 399.520 ;
        RECT 0.270 396.120 1377.175 396.760 ;
        RECT 4.400 394.720 1377.175 396.120 ;
        RECT 0.270 394.080 1377.175 394.720 ;
        RECT 4.400 391.320 1377.175 394.080 ;
        RECT 0.270 390.680 1377.175 391.320 ;
        RECT 4.400 389.280 1377.175 390.680 ;
        RECT 0.270 388.640 1377.175 389.280 ;
        RECT 4.400 385.880 1377.175 388.640 ;
        RECT 0.270 385.240 1377.175 385.880 ;
        RECT 4.400 382.480 1377.175 385.240 ;
        RECT 0.270 381.840 1377.175 382.480 ;
        RECT 4.400 380.440 1377.175 381.840 ;
        RECT 0.270 379.800 1377.175 380.440 ;
        RECT 4.400 377.040 1377.175 379.800 ;
        RECT 0.270 376.400 1377.175 377.040 ;
        RECT 4.400 375.000 1377.175 376.400 ;
        RECT 0.270 374.360 1377.175 375.000 ;
        RECT 4.400 371.600 1377.175 374.360 ;
        RECT 0.270 370.960 1377.175 371.600 ;
        RECT 4.400 369.560 1377.175 370.960 ;
        RECT 0.270 368.920 1377.175 369.560 ;
        RECT 4.400 366.160 1377.175 368.920 ;
        RECT 0.270 365.520 1377.175 366.160 ;
        RECT 4.400 362.760 1377.175 365.520 ;
        RECT 0.270 362.120 1377.175 362.760 ;
        RECT 4.400 360.720 1377.175 362.120 ;
        RECT 0.270 360.080 1377.175 360.720 ;
        RECT 4.400 357.320 1377.175 360.080 ;
        RECT 0.270 356.680 1377.175 357.320 ;
        RECT 4.400 355.280 1377.175 356.680 ;
        RECT 0.270 354.640 1377.175 355.280 ;
        RECT 4.400 351.880 1377.175 354.640 ;
        RECT 0.270 351.240 1377.175 351.880 ;
        RECT 4.400 348.480 1377.175 351.240 ;
        RECT 0.270 347.840 1377.175 348.480 ;
        RECT 4.400 346.440 1377.175 347.840 ;
        RECT 0.270 345.800 1377.175 346.440 ;
        RECT 4.400 343.040 1377.175 345.800 ;
        RECT 0.270 342.400 1377.175 343.040 ;
        RECT 4.400 341.000 1377.175 342.400 ;
        RECT 0.270 340.360 1377.175 341.000 ;
        RECT 4.400 337.600 1377.175 340.360 ;
        RECT 0.270 336.960 1377.175 337.600 ;
        RECT 4.400 334.200 1377.175 336.960 ;
        RECT 0.270 333.560 1377.175 334.200 ;
        RECT 4.400 332.160 1377.175 333.560 ;
        RECT 0.270 331.520 1377.175 332.160 ;
        RECT 4.400 328.760 1377.175 331.520 ;
        RECT 0.270 328.120 1377.175 328.760 ;
        RECT 4.400 326.720 1377.175 328.120 ;
        RECT 0.270 326.080 1377.175 326.720 ;
        RECT 4.400 323.320 1377.175 326.080 ;
        RECT 0.270 322.680 1377.175 323.320 ;
        RECT 4.400 319.920 1377.175 322.680 ;
        RECT 0.270 319.280 1377.175 319.920 ;
        RECT 4.400 317.880 1377.175 319.280 ;
        RECT 0.270 317.240 1377.175 317.880 ;
        RECT 4.400 314.480 1377.175 317.240 ;
        RECT 0.270 313.840 1377.175 314.480 ;
        RECT 4.400 312.440 1377.175 313.840 ;
        RECT 0.270 311.800 1377.175 312.440 ;
        RECT 4.400 309.040 1377.175 311.800 ;
        RECT 0.270 308.400 1377.175 309.040 ;
        RECT 4.400 305.640 1377.175 308.400 ;
        RECT 0.270 305.000 1377.175 305.640 ;
        RECT 4.400 303.600 1377.175 305.000 ;
        RECT 0.270 302.960 1377.175 303.600 ;
        RECT 4.400 300.200 1377.175 302.960 ;
        RECT 0.270 299.560 1377.175 300.200 ;
        RECT 4.400 298.160 1377.175 299.560 ;
        RECT 0.270 297.520 1377.175 298.160 ;
        RECT 4.400 294.760 1377.175 297.520 ;
        RECT 0.270 294.120 1377.175 294.760 ;
        RECT 4.400 291.360 1377.175 294.120 ;
        RECT 0.270 290.720 1377.175 291.360 ;
        RECT 4.400 289.320 1377.175 290.720 ;
        RECT 0.270 288.680 1377.175 289.320 ;
        RECT 4.400 285.920 1377.175 288.680 ;
        RECT 0.270 285.280 1377.175 285.920 ;
        RECT 4.400 283.880 1377.175 285.280 ;
        RECT 0.270 283.240 1377.175 283.880 ;
        RECT 4.400 280.480 1377.175 283.240 ;
        RECT 0.270 279.840 1377.175 280.480 ;
        RECT 4.400 277.080 1377.175 279.840 ;
        RECT 0.270 276.440 1377.175 277.080 ;
        RECT 4.400 275.040 1377.175 276.440 ;
        RECT 0.270 274.400 1377.175 275.040 ;
        RECT 4.400 271.640 1377.175 274.400 ;
        RECT 0.270 271.000 1377.175 271.640 ;
        RECT 4.400 269.600 1377.175 271.000 ;
        RECT 0.270 268.960 1377.175 269.600 ;
        RECT 4.400 266.200 1377.175 268.960 ;
        RECT 0.270 265.560 1377.175 266.200 ;
        RECT 4.400 262.800 1377.175 265.560 ;
        RECT 0.270 262.160 1377.175 262.800 ;
        RECT 4.400 260.760 1377.175 262.160 ;
        RECT 0.270 260.120 1377.175 260.760 ;
        RECT 4.400 257.360 1377.175 260.120 ;
        RECT 0.270 256.720 1377.175 257.360 ;
        RECT 4.400 255.320 1377.175 256.720 ;
        RECT 0.270 254.680 1377.175 255.320 ;
        RECT 4.400 251.920 1377.175 254.680 ;
        RECT 0.270 251.280 1377.175 251.920 ;
        RECT 4.400 248.520 1377.175 251.280 ;
        RECT 0.270 247.880 1377.175 248.520 ;
        RECT 4.400 246.480 1377.175 247.880 ;
        RECT 0.270 245.840 1377.175 246.480 ;
        RECT 4.400 243.080 1377.175 245.840 ;
        RECT 0.270 242.440 1377.175 243.080 ;
        RECT 4.400 241.040 1377.175 242.440 ;
        RECT 0.270 240.400 1377.175 241.040 ;
        RECT 4.400 237.640 1377.175 240.400 ;
        RECT 0.270 237.000 1377.175 237.640 ;
        RECT 4.400 234.240 1377.175 237.000 ;
        RECT 0.270 233.600 1377.175 234.240 ;
        RECT 4.400 232.200 1377.175 233.600 ;
        RECT 0.270 231.560 1377.175 232.200 ;
        RECT 4.400 228.800 1377.175 231.560 ;
        RECT 0.270 228.160 1377.175 228.800 ;
        RECT 4.400 226.760 1377.175 228.160 ;
        RECT 0.270 226.120 1377.175 226.760 ;
        RECT 4.400 223.360 1377.175 226.120 ;
        RECT 0.270 222.720 1377.175 223.360 ;
        RECT 4.400 219.960 1377.175 222.720 ;
        RECT 0.270 219.320 1377.175 219.960 ;
        RECT 4.400 217.920 1377.175 219.320 ;
        RECT 0.270 217.280 1377.175 217.920 ;
        RECT 4.400 214.520 1377.175 217.280 ;
        RECT 0.270 213.880 1377.175 214.520 ;
        RECT 4.400 212.480 1377.175 213.880 ;
        RECT 0.270 211.840 1377.175 212.480 ;
        RECT 4.400 209.080 1377.175 211.840 ;
        RECT 0.270 208.440 1377.175 209.080 ;
        RECT 4.400 205.680 1377.175 208.440 ;
        RECT 0.270 205.040 1377.175 205.680 ;
        RECT 4.400 203.640 1377.175 205.040 ;
        RECT 0.270 203.000 1377.175 203.640 ;
        RECT 4.400 200.240 1377.175 203.000 ;
        RECT 0.270 199.600 1377.175 200.240 ;
        RECT 4.400 198.200 1377.175 199.600 ;
        RECT 0.270 197.560 1377.175 198.200 ;
        RECT 4.400 194.800 1377.175 197.560 ;
        RECT 0.270 194.160 1377.175 194.800 ;
        RECT 4.400 191.400 1377.175 194.160 ;
        RECT 0.270 190.760 1377.175 191.400 ;
        RECT 4.400 189.360 1377.175 190.760 ;
        RECT 0.270 188.720 1377.175 189.360 ;
        RECT 4.400 185.960 1377.175 188.720 ;
        RECT 0.270 185.320 1377.175 185.960 ;
        RECT 4.400 183.920 1377.175 185.320 ;
        RECT 0.270 183.280 1377.175 183.920 ;
        RECT 4.400 180.520 1377.175 183.280 ;
        RECT 0.270 179.880 1377.175 180.520 ;
        RECT 4.400 178.480 1377.175 179.880 ;
        RECT 0.270 177.840 1377.175 178.480 ;
        RECT 4.400 175.080 1377.175 177.840 ;
        RECT 0.270 174.440 1377.175 175.080 ;
        RECT 4.400 171.680 1377.175 174.440 ;
        RECT 0.270 171.040 1377.175 171.680 ;
        RECT 4.400 169.640 1377.175 171.040 ;
        RECT 0.270 169.000 1377.175 169.640 ;
        RECT 4.400 166.240 1377.175 169.000 ;
        RECT 0.270 165.600 1377.175 166.240 ;
        RECT 4.400 164.200 1377.175 165.600 ;
        RECT 0.270 163.560 1377.175 164.200 ;
        RECT 4.400 160.800 1377.175 163.560 ;
        RECT 0.270 160.160 1377.175 160.800 ;
        RECT 4.400 157.400 1377.175 160.160 ;
        RECT 0.270 156.760 1377.175 157.400 ;
        RECT 4.400 155.360 1377.175 156.760 ;
        RECT 0.270 154.720 1377.175 155.360 ;
        RECT 4.400 151.960 1377.175 154.720 ;
        RECT 0.270 151.320 1377.175 151.960 ;
        RECT 4.400 149.920 1377.175 151.320 ;
        RECT 0.270 149.280 1377.175 149.920 ;
        RECT 4.400 146.520 1377.175 149.280 ;
        RECT 0.270 145.880 1377.175 146.520 ;
        RECT 4.400 143.120 1377.175 145.880 ;
        RECT 0.270 142.480 1377.175 143.120 ;
        RECT 4.400 141.080 1377.175 142.480 ;
        RECT 0.270 140.440 1377.175 141.080 ;
        RECT 4.400 137.680 1377.175 140.440 ;
        RECT 0.270 137.040 1377.175 137.680 ;
        RECT 4.400 135.640 1377.175 137.040 ;
        RECT 0.270 135.000 1377.175 135.640 ;
        RECT 4.400 132.240 1377.175 135.000 ;
        RECT 0.270 131.600 1377.175 132.240 ;
        RECT 4.400 128.840 1377.175 131.600 ;
        RECT 0.270 128.200 1377.175 128.840 ;
        RECT 4.400 126.800 1377.175 128.200 ;
        RECT 0.270 126.160 1377.175 126.800 ;
        RECT 4.400 123.400 1377.175 126.160 ;
        RECT 0.270 122.760 1377.175 123.400 ;
        RECT 4.400 121.360 1377.175 122.760 ;
        RECT 0.270 120.720 1377.175 121.360 ;
        RECT 4.400 117.960 1377.175 120.720 ;
        RECT 0.270 117.320 1377.175 117.960 ;
        RECT 4.400 114.560 1377.175 117.320 ;
        RECT 0.270 113.920 1377.175 114.560 ;
        RECT 4.400 112.520 1377.175 113.920 ;
        RECT 0.270 111.880 1377.175 112.520 ;
        RECT 4.400 109.120 1377.175 111.880 ;
        RECT 0.270 108.480 1377.175 109.120 ;
        RECT 4.400 107.080 1377.175 108.480 ;
        RECT 0.270 106.440 1377.175 107.080 ;
        RECT 4.400 103.680 1377.175 106.440 ;
        RECT 0.270 103.040 1377.175 103.680 ;
        RECT 4.400 100.280 1377.175 103.040 ;
        RECT 0.270 99.640 1377.175 100.280 ;
        RECT 4.400 98.240 1377.175 99.640 ;
        RECT 0.270 97.600 1377.175 98.240 ;
        RECT 4.400 94.840 1377.175 97.600 ;
        RECT 0.270 94.200 1377.175 94.840 ;
        RECT 4.400 92.800 1377.175 94.200 ;
        RECT 0.270 92.160 1377.175 92.800 ;
        RECT 4.400 89.400 1377.175 92.160 ;
        RECT 0.270 88.760 1377.175 89.400 ;
        RECT 4.400 86.000 1377.175 88.760 ;
        RECT 0.270 85.360 1377.175 86.000 ;
        RECT 4.400 83.960 1377.175 85.360 ;
        RECT 0.270 83.320 1377.175 83.960 ;
        RECT 4.400 80.560 1377.175 83.320 ;
        RECT 0.270 79.920 1377.175 80.560 ;
        RECT 4.400 78.520 1377.175 79.920 ;
        RECT 0.270 77.880 1377.175 78.520 ;
        RECT 4.400 75.120 1377.175 77.880 ;
        RECT 0.270 74.480 1377.175 75.120 ;
        RECT 4.400 71.720 1377.175 74.480 ;
        RECT 0.270 71.080 1377.175 71.720 ;
        RECT 4.400 69.680 1377.175 71.080 ;
        RECT 0.270 69.040 1377.175 69.680 ;
        RECT 4.400 66.280 1377.175 69.040 ;
        RECT 0.270 65.640 1377.175 66.280 ;
        RECT 4.400 64.240 1377.175 65.640 ;
        RECT 0.270 63.600 1377.175 64.240 ;
        RECT 4.400 60.840 1377.175 63.600 ;
        RECT 0.270 60.200 1377.175 60.840 ;
        RECT 4.400 57.440 1377.175 60.200 ;
        RECT 0.270 56.800 1377.175 57.440 ;
        RECT 4.400 55.400 1377.175 56.800 ;
        RECT 0.270 54.760 1377.175 55.400 ;
        RECT 4.400 52.000 1377.175 54.760 ;
        RECT 0.270 51.360 1377.175 52.000 ;
        RECT 4.400 49.960 1377.175 51.360 ;
        RECT 0.270 49.320 1377.175 49.960 ;
        RECT 4.400 46.560 1377.175 49.320 ;
        RECT 0.270 45.920 1377.175 46.560 ;
        RECT 4.400 43.160 1377.175 45.920 ;
        RECT 0.270 42.520 1377.175 43.160 ;
        RECT 4.400 41.120 1377.175 42.520 ;
        RECT 0.270 40.480 1377.175 41.120 ;
        RECT 4.400 37.720 1377.175 40.480 ;
        RECT 0.270 37.080 1377.175 37.720 ;
        RECT 4.400 35.680 1377.175 37.080 ;
        RECT 0.270 35.040 1377.175 35.680 ;
        RECT 4.400 32.280 1377.175 35.040 ;
        RECT 0.270 31.640 1377.175 32.280 ;
        RECT 4.400 28.880 1377.175 31.640 ;
        RECT 0.270 28.240 1377.175 28.880 ;
        RECT 4.400 26.840 1377.175 28.240 ;
        RECT 0.270 26.200 1377.175 26.840 ;
        RECT 4.400 23.440 1377.175 26.200 ;
        RECT 0.270 22.800 1377.175 23.440 ;
        RECT 4.400 21.400 1377.175 22.800 ;
        RECT 0.270 20.760 1377.175 21.400 ;
        RECT 4.400 18.000 1377.175 20.760 ;
        RECT 0.270 17.360 1377.175 18.000 ;
        RECT 4.400 14.600 1377.175 17.360 ;
        RECT 0.270 13.960 1377.175 14.600 ;
        RECT 4.400 12.560 1377.175 13.960 ;
        RECT 0.270 11.920 1377.175 12.560 ;
        RECT 4.400 9.160 1377.175 11.920 ;
        RECT 0.270 8.520 1377.175 9.160 ;
        RECT 4.400 7.120 1377.175 8.520 ;
        RECT 0.270 6.480 1377.175 7.120 ;
        RECT 4.400 3.720 1377.175 6.480 ;
        RECT 0.270 3.080 1377.175 3.720 ;
        RECT 4.400 0.855 1377.175 3.080 ;
      LAYER met4 ;
        RECT 0.295 1488.480 1367.745 1497.185 ;
        RECT 0.295 10.240 20.640 1488.480 ;
        RECT 23.040 10.240 97.440 1488.480 ;
        RECT 99.840 10.240 174.240 1488.480 ;
        RECT 176.640 10.240 251.040 1488.480 ;
        RECT 253.440 10.240 327.840 1488.480 ;
        RECT 330.240 10.240 404.640 1488.480 ;
        RECT 407.040 10.240 481.440 1488.480 ;
        RECT 483.840 10.240 558.240 1488.480 ;
        RECT 560.640 10.240 635.040 1488.480 ;
        RECT 637.440 10.240 711.840 1488.480 ;
        RECT 714.240 10.240 788.640 1488.480 ;
        RECT 791.040 10.240 865.440 1488.480 ;
        RECT 867.840 10.240 942.240 1488.480 ;
        RECT 944.640 10.240 1019.040 1488.480 ;
        RECT 1021.440 10.240 1095.840 1488.480 ;
        RECT 1098.240 10.240 1172.640 1488.480 ;
        RECT 1175.040 10.240 1249.440 1488.480 ;
        RECT 1251.840 10.240 1326.240 1488.480 ;
        RECT 1328.640 10.240 1367.745 1488.480 ;
        RECT 0.295 9.015 1367.745 10.240 ;
  END
END el2_swerv_wrapper
END LIBRARY

