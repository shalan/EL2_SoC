magic
tech sky130A
magscale 1 2
timestamp 1611159231
<< obsli1 >>
rect 442 2159 158377 157777
<< obsm1 >>
rect 442 1436 158576 157808
<< metal2 >>
rect 0 159200 56 160000
rect 1380 159200 1436 160000
rect 2852 159200 2908 160000
rect 4232 159200 4288 160000
rect 5704 159200 5760 160000
rect 7084 159200 7140 160000
rect 8556 159200 8612 160000
rect 9936 159200 9992 160000
rect 11408 159200 11464 160000
rect 12788 159200 12844 160000
rect 14260 159200 14316 160000
rect 15640 159200 15696 160000
rect 17112 159200 17168 160000
rect 18492 159200 18548 160000
rect 19964 159200 20020 160000
rect 21344 159200 21400 160000
rect 22816 159200 22872 160000
rect 24196 159200 24252 160000
rect 25668 159200 25724 160000
rect 27140 159200 27196 160000
rect 28520 159200 28576 160000
rect 29992 159200 30048 160000
rect 31372 159200 31428 160000
rect 32844 159200 32900 160000
rect 34224 159200 34280 160000
rect 35696 159200 35752 160000
rect 37076 159200 37132 160000
rect 38548 159200 38604 160000
rect 39928 159200 39984 160000
rect 41400 159200 41456 160000
rect 42780 159200 42836 160000
rect 44252 159200 44308 160000
rect 45632 159200 45688 160000
rect 47104 159200 47160 160000
rect 48484 159200 48540 160000
rect 49956 159200 50012 160000
rect 51336 159200 51392 160000
rect 52808 159200 52864 160000
rect 54280 159200 54336 160000
rect 55660 159200 55716 160000
rect 57132 159200 57188 160000
rect 58512 159200 58568 160000
rect 59984 159200 60040 160000
rect 61364 159200 61420 160000
rect 62836 159200 62892 160000
rect 64216 159200 64272 160000
rect 65688 159200 65744 160000
rect 67068 159200 67124 160000
rect 68540 159200 68596 160000
rect 69920 159200 69976 160000
rect 71392 159200 71448 160000
rect 72772 159200 72828 160000
rect 74244 159200 74300 160000
rect 75624 159200 75680 160000
rect 77096 159200 77152 160000
rect 78476 159200 78532 160000
rect 79948 159200 80004 160000
rect 81420 159200 81476 160000
rect 82800 159200 82856 160000
rect 84272 159200 84328 160000
rect 85652 159200 85708 160000
rect 87124 159200 87180 160000
rect 88504 159200 88560 160000
rect 89976 159200 90032 160000
rect 91356 159200 91412 160000
rect 92828 159200 92884 160000
rect 94208 159200 94264 160000
rect 95680 159200 95736 160000
rect 97060 159200 97116 160000
rect 98532 159200 98588 160000
rect 99912 159200 99968 160000
rect 101384 159200 101440 160000
rect 102764 159200 102820 160000
rect 104236 159200 104292 160000
rect 105616 159200 105672 160000
rect 107088 159200 107144 160000
rect 108560 159200 108616 160000
rect 109940 159200 109996 160000
rect 111412 159200 111468 160000
rect 112792 159200 112848 160000
rect 114264 159200 114320 160000
rect 115644 159200 115700 160000
rect 117116 159200 117172 160000
rect 118496 159200 118552 160000
rect 119968 159200 120024 160000
rect 121348 159200 121404 160000
rect 122820 159200 122876 160000
rect 124200 159200 124256 160000
rect 125672 159200 125728 160000
rect 127052 159200 127108 160000
rect 128524 159200 128580 160000
rect 129904 159200 129960 160000
rect 131376 159200 131432 160000
rect 132756 159200 132812 160000
rect 134228 159200 134284 160000
rect 135700 159200 135756 160000
rect 137080 159200 137136 160000
rect 138552 159200 138608 160000
rect 139932 159200 139988 160000
rect 141404 159200 141460 160000
rect 142784 159200 142840 160000
rect 144256 159200 144312 160000
rect 145636 159200 145692 160000
rect 147108 159200 147164 160000
rect 148488 159200 148544 160000
rect 149960 159200 150016 160000
rect 151340 159200 151396 160000
rect 152812 159200 152868 160000
rect 154192 159200 154248 160000
rect 155664 159200 155720 160000
rect 157044 159200 157100 160000
rect 158516 159200 158572 160000
rect 19320 0 19376 800
rect 59248 0 59304 800
rect 99268 0 99324 800
rect 139288 0 139344 800
<< obsm2 >>
rect 3558 159144 4176 159225
rect 4344 159144 5648 159225
rect 5816 159144 7028 159225
rect 7196 159144 8500 159225
rect 8668 159144 9880 159225
rect 10048 159144 11352 159225
rect 11520 159144 12732 159225
rect 12900 159144 14204 159225
rect 14372 159144 15584 159225
rect 15752 159144 17056 159225
rect 17224 159144 18436 159225
rect 18604 159144 19908 159225
rect 20076 159144 21288 159225
rect 21456 159144 22760 159225
rect 22928 159144 24140 159225
rect 24308 159144 25612 159225
rect 25780 159144 27084 159225
rect 27252 159144 28464 159225
rect 28632 159144 29936 159225
rect 30104 159144 31316 159225
rect 31484 159144 32788 159225
rect 32956 159144 34168 159225
rect 34336 159144 35640 159225
rect 35808 159144 37020 159225
rect 37188 159144 38492 159225
rect 38660 159144 39872 159225
rect 40040 159144 41344 159225
rect 41512 159144 42724 159225
rect 42892 159144 44196 159225
rect 44364 159144 45576 159225
rect 45744 159144 47048 159225
rect 47216 159144 48428 159225
rect 48596 159144 49900 159225
rect 50068 159144 51280 159225
rect 51448 159144 52752 159225
rect 52920 159144 54224 159225
rect 54392 159144 55604 159225
rect 55772 159144 57076 159225
rect 57244 159144 58456 159225
rect 58624 159144 59928 159225
rect 60096 159144 61308 159225
rect 61476 159144 62780 159225
rect 62948 159144 64160 159225
rect 64328 159144 65632 159225
rect 65800 159144 67012 159225
rect 67180 159144 68484 159225
rect 68652 159144 69864 159225
rect 70032 159144 71336 159225
rect 71504 159144 72716 159225
rect 72884 159144 74188 159225
rect 74356 159144 75568 159225
rect 75736 159144 77040 159225
rect 77208 159144 78420 159225
rect 78588 159144 79892 159225
rect 80060 159144 81364 159225
rect 81532 159144 82744 159225
rect 82912 159144 84216 159225
rect 84384 159144 85596 159225
rect 85764 159144 87068 159225
rect 87236 159144 88448 159225
rect 88616 159144 89920 159225
rect 90088 159144 91300 159225
rect 91468 159144 92772 159225
rect 92940 159144 94152 159225
rect 94320 159144 95624 159225
rect 95792 159144 97004 159225
rect 97172 159144 98476 159225
rect 98644 159144 99856 159225
rect 100024 159144 101328 159225
rect 101496 159144 102708 159225
rect 102876 159144 104180 159225
rect 104348 159144 105560 159225
rect 105728 159144 107032 159225
rect 107200 159144 108504 159225
rect 108672 159144 109884 159225
rect 110052 159144 111356 159225
rect 111524 159144 112736 159225
rect 112904 159144 114208 159225
rect 114376 159144 115588 159225
rect 115756 159144 117060 159225
rect 117228 159144 118440 159225
rect 118608 159144 119912 159225
rect 120080 159144 121292 159225
rect 121460 159144 122764 159225
rect 122932 159144 124144 159225
rect 124312 159144 125616 159225
rect 125784 159144 126996 159225
rect 127164 159144 128468 159225
rect 128636 159144 129848 159225
rect 130016 159144 131320 159225
rect 131488 159144 132700 159225
rect 132868 159144 134172 159225
rect 134340 159144 135644 159225
rect 135812 159144 137024 159225
rect 137192 159144 138496 159225
rect 138664 159144 139876 159225
rect 140044 159144 141348 159225
rect 141516 159144 142728 159225
rect 142896 159144 144200 159225
rect 144368 159144 145580 159225
rect 145748 159144 147052 159225
rect 147220 159144 148432 159225
rect 148600 159144 149904 159225
rect 150072 159144 151284 159225
rect 151452 159144 152756 159225
rect 152924 159144 154136 159225
rect 154304 159144 155608 159225
rect 155776 159144 156988 159225
rect 157156 159144 158460 159225
rect 3558 856 158570 159144
rect 3558 800 19264 856
rect 19432 800 59192 856
rect 59360 800 99212 856
rect 99380 800 139232 856
rect 139400 800 158570 856
<< metal3 >>
rect 158538 159128 159338 159248
rect 158538 157904 159338 158024
rect 158538 156680 159338 156800
rect 158538 155456 159338 155576
rect 158538 154232 159338 154352
rect 158538 152872 159338 152992
rect 158538 151648 159338 151768
rect 158538 150424 159338 150544
rect 158538 149200 159338 149320
rect 158538 147976 159338 148096
rect 158538 146616 159338 146736
rect 158538 145392 159338 145512
rect 158538 144168 159338 144288
rect 158538 142944 159338 143064
rect 158538 141720 159338 141840
rect 158538 140496 159338 140616
rect 158538 139136 159338 139256
rect 158538 137912 159338 138032
rect 158538 136688 159338 136808
rect 158538 135464 159338 135584
rect 158538 134240 159338 134360
rect 158538 132880 159338 133000
rect 158538 131656 159338 131776
rect 158538 130432 159338 130552
rect 158538 129208 159338 129328
rect 158538 127984 159338 128104
rect 158538 126624 159338 126744
rect 158538 125400 159338 125520
rect 158538 124176 159338 124296
rect 158538 122952 159338 123072
rect 158538 121728 159338 121848
rect 158538 120504 159338 120624
rect 158538 119144 159338 119264
rect 158538 117920 159338 118040
rect 158538 116696 159338 116816
rect 158538 115472 159338 115592
rect 158538 114248 159338 114368
rect 158538 112888 159338 113008
rect 158538 111664 159338 111784
rect 158538 110440 159338 110560
rect 158538 109216 159338 109336
rect 158538 107992 159338 108112
rect 158538 106632 159338 106752
rect 158538 105408 159338 105528
rect 158538 104184 159338 104304
rect 158538 102960 159338 103080
rect 158538 101736 159338 101856
rect 158538 100512 159338 100632
rect 158538 99152 159338 99272
rect 158538 97928 159338 98048
rect 158538 96704 159338 96824
rect 158538 95480 159338 95600
rect 158538 94256 159338 94376
rect 158538 92896 159338 93016
rect 158538 91672 159338 91792
rect 158538 90448 159338 90568
rect 158538 89224 159338 89344
rect 158538 88000 159338 88120
rect 158538 86640 159338 86760
rect 158538 85416 159338 85536
rect 158538 84192 159338 84312
rect 158538 82968 159338 83088
rect 158538 81744 159338 81864
rect 158538 80520 159338 80640
rect 158538 79160 159338 79280
rect 158538 77936 159338 78056
rect 158538 76712 159338 76832
rect 158538 75488 159338 75608
rect 158538 74264 159338 74384
rect 158538 72904 159338 73024
rect 158538 71680 159338 71800
rect 158538 70456 159338 70576
rect 158538 69232 159338 69352
rect 158538 68008 159338 68128
rect 158538 66648 159338 66768
rect 158538 65424 159338 65544
rect 158538 64200 159338 64320
rect 158538 62976 159338 63096
rect 158538 61752 159338 61872
rect 158538 60528 159338 60648
rect 158538 59168 159338 59288
rect 158538 57944 159338 58064
rect 158538 56720 159338 56840
rect 158538 55496 159338 55616
rect 158538 54272 159338 54392
rect 158538 52912 159338 53032
rect 158538 51688 159338 51808
rect 158538 50464 159338 50584
rect 158538 49240 159338 49360
rect 158538 48016 159338 48136
rect 158538 46656 159338 46776
rect 158538 45432 159338 45552
rect 158538 44208 159338 44328
rect 158538 42984 159338 43104
rect 158538 41760 159338 41880
rect 158538 40536 159338 40656
rect 158538 39176 159338 39296
rect 158538 37952 159338 38072
rect 158538 36728 159338 36848
rect 158538 35504 159338 35624
rect 158538 34280 159338 34400
rect 158538 32920 159338 33040
rect 158538 31696 159338 31816
rect 158538 30472 159338 30592
rect 158538 29248 159338 29368
rect 158538 28024 159338 28144
rect 158538 26664 159338 26784
rect 158538 25440 159338 25560
rect 158538 24216 159338 24336
rect 158538 22992 159338 23112
rect 158538 21768 159338 21888
rect 158538 20544 159338 20664
rect 158538 19184 159338 19304
rect 158538 17960 159338 18080
rect 158538 16736 159338 16856
rect 158538 15512 159338 15632
rect 158538 14288 159338 14408
rect 158538 12928 159338 13048
rect 158538 11704 159338 11824
rect 158538 10480 159338 10600
rect 158538 9256 159338 9376
rect 158538 8032 159338 8152
rect 158538 6672 159338 6792
rect 158538 5448 159338 5568
rect 158538 4224 159338 4344
rect 158538 3000 159338 3120
rect 158538 1776 159338 1896
rect 158538 552 159338 672
<< obsm3 >>
rect 3546 159048 158458 159221
rect 3546 158104 158538 159048
rect 3546 157824 158458 158104
rect 3546 156880 158538 157824
rect 3546 156600 158458 156880
rect 3546 155656 158538 156600
rect 3546 155376 158458 155656
rect 3546 154432 158538 155376
rect 3546 154152 158458 154432
rect 3546 153072 158538 154152
rect 3546 152792 158458 153072
rect 3546 151848 158538 152792
rect 3546 151568 158458 151848
rect 3546 150624 158538 151568
rect 3546 150344 158458 150624
rect 3546 149400 158538 150344
rect 3546 149120 158458 149400
rect 3546 148176 158538 149120
rect 3546 147896 158458 148176
rect 3546 146816 158538 147896
rect 3546 146536 158458 146816
rect 3546 145592 158538 146536
rect 3546 145312 158458 145592
rect 3546 144368 158538 145312
rect 3546 144088 158458 144368
rect 3546 143144 158538 144088
rect 3546 142864 158458 143144
rect 3546 141920 158538 142864
rect 3546 141640 158458 141920
rect 3546 140696 158538 141640
rect 3546 140416 158458 140696
rect 3546 139336 158538 140416
rect 3546 139056 158458 139336
rect 3546 138112 158538 139056
rect 3546 137832 158458 138112
rect 3546 136888 158538 137832
rect 3546 136608 158458 136888
rect 3546 135664 158538 136608
rect 3546 135384 158458 135664
rect 3546 134440 158538 135384
rect 3546 134160 158458 134440
rect 3546 133080 158538 134160
rect 3546 132800 158458 133080
rect 3546 131856 158538 132800
rect 3546 131576 158458 131856
rect 3546 130632 158538 131576
rect 3546 130352 158458 130632
rect 3546 129408 158538 130352
rect 3546 129128 158458 129408
rect 3546 128184 158538 129128
rect 3546 127904 158458 128184
rect 3546 126824 158538 127904
rect 3546 126544 158458 126824
rect 3546 125600 158538 126544
rect 3546 125320 158458 125600
rect 3546 124376 158538 125320
rect 3546 124096 158458 124376
rect 3546 123152 158538 124096
rect 3546 122872 158458 123152
rect 3546 121928 158538 122872
rect 3546 121648 158458 121928
rect 3546 120704 158538 121648
rect 3546 120424 158458 120704
rect 3546 119344 158538 120424
rect 3546 119064 158458 119344
rect 3546 118120 158538 119064
rect 3546 117840 158458 118120
rect 3546 116896 158538 117840
rect 3546 116616 158458 116896
rect 3546 115672 158538 116616
rect 3546 115392 158458 115672
rect 3546 114448 158538 115392
rect 3546 114168 158458 114448
rect 3546 113088 158538 114168
rect 3546 112808 158458 113088
rect 3546 111864 158538 112808
rect 3546 111584 158458 111864
rect 3546 110640 158538 111584
rect 3546 110360 158458 110640
rect 3546 109416 158538 110360
rect 3546 109136 158458 109416
rect 3546 108192 158538 109136
rect 3546 107912 158458 108192
rect 3546 106832 158538 107912
rect 3546 106552 158458 106832
rect 3546 105608 158538 106552
rect 3546 105328 158458 105608
rect 3546 104384 158538 105328
rect 3546 104104 158458 104384
rect 3546 103160 158538 104104
rect 3546 102880 158458 103160
rect 3546 101936 158538 102880
rect 3546 101656 158458 101936
rect 3546 100712 158538 101656
rect 3546 100432 158458 100712
rect 3546 99352 158538 100432
rect 3546 99072 158458 99352
rect 3546 98128 158538 99072
rect 3546 97848 158458 98128
rect 3546 96904 158538 97848
rect 3546 96624 158458 96904
rect 3546 95680 158538 96624
rect 3546 95400 158458 95680
rect 3546 94456 158538 95400
rect 3546 94176 158458 94456
rect 3546 93096 158538 94176
rect 3546 92816 158458 93096
rect 3546 91872 158538 92816
rect 3546 91592 158458 91872
rect 3546 90648 158538 91592
rect 3546 90368 158458 90648
rect 3546 89424 158538 90368
rect 3546 89144 158458 89424
rect 3546 88200 158538 89144
rect 3546 87920 158458 88200
rect 3546 86840 158538 87920
rect 3546 86560 158458 86840
rect 3546 85616 158538 86560
rect 3546 85336 158458 85616
rect 3546 84392 158538 85336
rect 3546 84112 158458 84392
rect 3546 83168 158538 84112
rect 3546 82888 158458 83168
rect 3546 81944 158538 82888
rect 3546 81664 158458 81944
rect 3546 80720 158538 81664
rect 3546 80440 158458 80720
rect 3546 79360 158538 80440
rect 3546 79080 158458 79360
rect 3546 78136 158538 79080
rect 3546 77856 158458 78136
rect 3546 76912 158538 77856
rect 3546 76632 158458 76912
rect 3546 75688 158538 76632
rect 3546 75408 158458 75688
rect 3546 74464 158538 75408
rect 3546 74184 158458 74464
rect 3546 73104 158538 74184
rect 3546 72824 158458 73104
rect 3546 71880 158538 72824
rect 3546 71600 158458 71880
rect 3546 70656 158538 71600
rect 3546 70376 158458 70656
rect 3546 69432 158538 70376
rect 3546 69152 158458 69432
rect 3546 68208 158538 69152
rect 3546 67928 158458 68208
rect 3546 66848 158538 67928
rect 3546 66568 158458 66848
rect 3546 65624 158538 66568
rect 3546 65344 158458 65624
rect 3546 64400 158538 65344
rect 3546 64120 158458 64400
rect 3546 63176 158538 64120
rect 3546 62896 158458 63176
rect 3546 61952 158538 62896
rect 3546 61672 158458 61952
rect 3546 60728 158538 61672
rect 3546 60448 158458 60728
rect 3546 59368 158538 60448
rect 3546 59088 158458 59368
rect 3546 58144 158538 59088
rect 3546 57864 158458 58144
rect 3546 56920 158538 57864
rect 3546 56640 158458 56920
rect 3546 55696 158538 56640
rect 3546 55416 158458 55696
rect 3546 54472 158538 55416
rect 3546 54192 158458 54472
rect 3546 53112 158538 54192
rect 3546 52832 158458 53112
rect 3546 51888 158538 52832
rect 3546 51608 158458 51888
rect 3546 50664 158538 51608
rect 3546 50384 158458 50664
rect 3546 49440 158538 50384
rect 3546 49160 158458 49440
rect 3546 48216 158538 49160
rect 3546 47936 158458 48216
rect 3546 46856 158538 47936
rect 3546 46576 158458 46856
rect 3546 45632 158538 46576
rect 3546 45352 158458 45632
rect 3546 44408 158538 45352
rect 3546 44128 158458 44408
rect 3546 43184 158538 44128
rect 3546 42904 158458 43184
rect 3546 41960 158538 42904
rect 3546 41680 158458 41960
rect 3546 40736 158538 41680
rect 3546 40456 158458 40736
rect 3546 39376 158538 40456
rect 3546 39096 158458 39376
rect 3546 38152 158538 39096
rect 3546 37872 158458 38152
rect 3546 36928 158538 37872
rect 3546 36648 158458 36928
rect 3546 35704 158538 36648
rect 3546 35424 158458 35704
rect 3546 34480 158538 35424
rect 3546 34200 158458 34480
rect 3546 33120 158538 34200
rect 3546 32840 158458 33120
rect 3546 31896 158538 32840
rect 3546 31616 158458 31896
rect 3546 30672 158538 31616
rect 3546 30392 158458 30672
rect 3546 29448 158538 30392
rect 3546 29168 158458 29448
rect 3546 28224 158538 29168
rect 3546 27944 158458 28224
rect 3546 26864 158538 27944
rect 3546 26584 158458 26864
rect 3546 25640 158538 26584
rect 3546 25360 158458 25640
rect 3546 24416 158538 25360
rect 3546 24136 158458 24416
rect 3546 23192 158538 24136
rect 3546 22912 158458 23192
rect 3546 21968 158538 22912
rect 3546 21688 158458 21968
rect 3546 20744 158538 21688
rect 3546 20464 158458 20744
rect 3546 19384 158538 20464
rect 3546 19104 158458 19384
rect 3546 18160 158538 19104
rect 3546 17880 158458 18160
rect 3546 16936 158538 17880
rect 3546 16656 158458 16936
rect 3546 15712 158538 16656
rect 3546 15432 158458 15712
rect 3546 14488 158538 15432
rect 3546 14208 158458 14488
rect 3546 13128 158538 14208
rect 3546 12848 158458 13128
rect 3546 11904 158538 12848
rect 3546 11624 158458 11904
rect 3546 10680 158538 11624
rect 3546 10400 158458 10680
rect 3546 9456 158538 10400
rect 3546 9176 158458 9456
rect 3546 8232 158538 9176
rect 3546 7952 158458 8232
rect 3546 6872 158538 7952
rect 3546 6592 158458 6872
rect 3546 5648 158538 6592
rect 3546 5368 158458 5648
rect 3546 4424 158538 5368
rect 3546 4144 158458 4424
rect 3546 3200 158538 4144
rect 3546 2920 158458 3200
rect 3546 1976 158538 2920
rect 3546 1696 158458 1976
rect 3546 752 158538 1696
rect 3546 472 158458 752
rect 3546 36 158538 472
<< metal4 >>
rect 3546 2128 3866 157808
rect 18906 2128 19226 157808
rect 34266 2128 34586 157808
rect 49626 2128 49946 157808
rect 64986 2128 65306 157808
rect 80346 2128 80666 157808
rect 95706 2128 96026 157808
rect 111066 2128 111386 157808
rect 126426 2128 126746 157808
rect 141786 2128 142106 157808
rect 157146 2128 157466 157808
<< obsm4 >>
rect 27365 2048 34186 157589
rect 34666 2048 49546 157589
rect 50026 2048 64906 157589
rect 65386 2048 80266 157589
rect 80746 2048 95626 157589
rect 96106 2048 110986 157589
rect 111466 2048 126346 157589
rect 126826 2048 141706 157589
rect 142186 2048 155127 157589
rect 27365 35 155127 2048
<< labels >>
rlabel metal2 s 0 159200 56 160000 6 A[0]
port 1 nsew signal input
rlabel metal2 s 14260 159200 14316 160000 6 A[10]
port 2 nsew signal input
rlabel metal2 s 15640 159200 15696 160000 6 A[11]
port 3 nsew signal input
rlabel metal2 s 17112 159200 17168 160000 6 A[12]
port 4 nsew signal input
rlabel metal2 s 18492 159200 18548 160000 6 A[13]
port 5 nsew signal input
rlabel metal2 s 19964 159200 20020 160000 6 A[14]
port 6 nsew signal input
rlabel metal2 s 21344 159200 21400 160000 6 A[15]
port 7 nsew signal input
rlabel metal2 s 22816 159200 22872 160000 6 A[16]
port 8 nsew signal input
rlabel metal2 s 24196 159200 24252 160000 6 A[17]
port 9 nsew signal input
rlabel metal2 s 25668 159200 25724 160000 6 A[18]
port 10 nsew signal input
rlabel metal2 s 27140 159200 27196 160000 6 A[19]
port 11 nsew signal input
rlabel metal2 s 1380 159200 1436 160000 6 A[1]
port 12 nsew signal input
rlabel metal2 s 28520 159200 28576 160000 6 A[20]
port 13 nsew signal input
rlabel metal2 s 29992 159200 30048 160000 6 A[21]
port 14 nsew signal input
rlabel metal2 s 31372 159200 31428 160000 6 A[22]
port 15 nsew signal input
rlabel metal2 s 32844 159200 32900 160000 6 A[23]
port 16 nsew signal input
rlabel metal2 s 2852 159200 2908 160000 6 A[2]
port 17 nsew signal input
rlabel metal2 s 4232 159200 4288 160000 6 A[3]
port 18 nsew signal input
rlabel metal2 s 5704 159200 5760 160000 6 A[4]
port 19 nsew signal input
rlabel metal2 s 7084 159200 7140 160000 6 A[5]
port 20 nsew signal input
rlabel metal2 s 8556 159200 8612 160000 6 A[6]
port 21 nsew signal input
rlabel metal2 s 9936 159200 9992 160000 6 A[7]
port 22 nsew signal input
rlabel metal2 s 11408 159200 11464 160000 6 A[8]
port 23 nsew signal input
rlabel metal2 s 12788 159200 12844 160000 6 A[9]
port 24 nsew signal input
rlabel metal2 s 34224 159200 34280 160000 6 A_h[0]
port 25 nsew signal input
rlabel metal2 s 48484 159200 48540 160000 6 A_h[10]
port 26 nsew signal input
rlabel metal2 s 49956 159200 50012 160000 6 A_h[11]
port 27 nsew signal input
rlabel metal2 s 51336 159200 51392 160000 6 A_h[12]
port 28 nsew signal input
rlabel metal2 s 52808 159200 52864 160000 6 A_h[13]
port 29 nsew signal input
rlabel metal2 s 54280 159200 54336 160000 6 A_h[14]
port 30 nsew signal input
rlabel metal2 s 55660 159200 55716 160000 6 A_h[15]
port 31 nsew signal input
rlabel metal2 s 57132 159200 57188 160000 6 A_h[16]
port 32 nsew signal input
rlabel metal2 s 58512 159200 58568 160000 6 A_h[17]
port 33 nsew signal input
rlabel metal2 s 59984 159200 60040 160000 6 A_h[18]
port 34 nsew signal input
rlabel metal2 s 61364 159200 61420 160000 6 A_h[19]
port 35 nsew signal input
rlabel metal2 s 35696 159200 35752 160000 6 A_h[1]
port 36 nsew signal input
rlabel metal2 s 62836 159200 62892 160000 6 A_h[20]
port 37 nsew signal input
rlabel metal2 s 64216 159200 64272 160000 6 A_h[21]
port 38 nsew signal input
rlabel metal2 s 65688 159200 65744 160000 6 A_h[22]
port 39 nsew signal input
rlabel metal2 s 67068 159200 67124 160000 6 A_h[23]
port 40 nsew signal input
rlabel metal2 s 37076 159200 37132 160000 6 A_h[2]
port 41 nsew signal input
rlabel metal2 s 38548 159200 38604 160000 6 A_h[3]
port 42 nsew signal input
rlabel metal2 s 39928 159200 39984 160000 6 A_h[4]
port 43 nsew signal input
rlabel metal2 s 41400 159200 41456 160000 6 A_h[5]
port 44 nsew signal input
rlabel metal2 s 42780 159200 42836 160000 6 A_h[6]
port 45 nsew signal input
rlabel metal2 s 44252 159200 44308 160000 6 A_h[7]
port 46 nsew signal input
rlabel metal2 s 45632 159200 45688 160000 6 A_h[8]
port 47 nsew signal input
rlabel metal2 s 47104 159200 47160 160000 6 A_h[9]
port 48 nsew signal input
rlabel metal2 s 68540 159200 68596 160000 6 Do[0]
port 49 nsew signal output
rlabel metal2 s 82800 159200 82856 160000 6 Do[10]
port 50 nsew signal output
rlabel metal2 s 84272 159200 84328 160000 6 Do[11]
port 51 nsew signal output
rlabel metal2 s 85652 159200 85708 160000 6 Do[12]
port 52 nsew signal output
rlabel metal2 s 87124 159200 87180 160000 6 Do[13]
port 53 nsew signal output
rlabel metal2 s 88504 159200 88560 160000 6 Do[14]
port 54 nsew signal output
rlabel metal2 s 89976 159200 90032 160000 6 Do[15]
port 55 nsew signal output
rlabel metal2 s 91356 159200 91412 160000 6 Do[16]
port 56 nsew signal output
rlabel metal2 s 92828 159200 92884 160000 6 Do[17]
port 57 nsew signal output
rlabel metal2 s 94208 159200 94264 160000 6 Do[18]
port 58 nsew signal output
rlabel metal2 s 95680 159200 95736 160000 6 Do[19]
port 59 nsew signal output
rlabel metal2 s 69920 159200 69976 160000 6 Do[1]
port 60 nsew signal output
rlabel metal2 s 97060 159200 97116 160000 6 Do[20]
port 61 nsew signal output
rlabel metal2 s 98532 159200 98588 160000 6 Do[21]
port 62 nsew signal output
rlabel metal2 s 99912 159200 99968 160000 6 Do[22]
port 63 nsew signal output
rlabel metal2 s 101384 159200 101440 160000 6 Do[23]
port 64 nsew signal output
rlabel metal2 s 102764 159200 102820 160000 6 Do[24]
port 65 nsew signal output
rlabel metal2 s 104236 159200 104292 160000 6 Do[25]
port 66 nsew signal output
rlabel metal2 s 105616 159200 105672 160000 6 Do[26]
port 67 nsew signal output
rlabel metal2 s 107088 159200 107144 160000 6 Do[27]
port 68 nsew signal output
rlabel metal2 s 108560 159200 108616 160000 6 Do[28]
port 69 nsew signal output
rlabel metal2 s 109940 159200 109996 160000 6 Do[29]
port 70 nsew signal output
rlabel metal2 s 71392 159200 71448 160000 6 Do[2]
port 71 nsew signal output
rlabel metal2 s 111412 159200 111468 160000 6 Do[30]
port 72 nsew signal output
rlabel metal2 s 112792 159200 112848 160000 6 Do[31]
port 73 nsew signal output
rlabel metal2 s 114264 159200 114320 160000 6 Do[32]
port 74 nsew signal output
rlabel metal2 s 115644 159200 115700 160000 6 Do[33]
port 75 nsew signal output
rlabel metal2 s 117116 159200 117172 160000 6 Do[34]
port 76 nsew signal output
rlabel metal2 s 118496 159200 118552 160000 6 Do[35]
port 77 nsew signal output
rlabel metal2 s 119968 159200 120024 160000 6 Do[36]
port 78 nsew signal output
rlabel metal2 s 121348 159200 121404 160000 6 Do[37]
port 79 nsew signal output
rlabel metal2 s 122820 159200 122876 160000 6 Do[38]
port 80 nsew signal output
rlabel metal2 s 124200 159200 124256 160000 6 Do[39]
port 81 nsew signal output
rlabel metal2 s 72772 159200 72828 160000 6 Do[3]
port 82 nsew signal output
rlabel metal2 s 125672 159200 125728 160000 6 Do[40]
port 83 nsew signal output
rlabel metal2 s 127052 159200 127108 160000 6 Do[41]
port 84 nsew signal output
rlabel metal2 s 128524 159200 128580 160000 6 Do[42]
port 85 nsew signal output
rlabel metal2 s 129904 159200 129960 160000 6 Do[43]
port 86 nsew signal output
rlabel metal2 s 131376 159200 131432 160000 6 Do[44]
port 87 nsew signal output
rlabel metal2 s 132756 159200 132812 160000 6 Do[45]
port 88 nsew signal output
rlabel metal2 s 134228 159200 134284 160000 6 Do[46]
port 89 nsew signal output
rlabel metal2 s 135700 159200 135756 160000 6 Do[47]
port 90 nsew signal output
rlabel metal2 s 137080 159200 137136 160000 6 Do[48]
port 91 nsew signal output
rlabel metal2 s 138552 159200 138608 160000 6 Do[49]
port 92 nsew signal output
rlabel metal2 s 74244 159200 74300 160000 6 Do[4]
port 93 nsew signal output
rlabel metal2 s 139932 159200 139988 160000 6 Do[50]
port 94 nsew signal output
rlabel metal2 s 141404 159200 141460 160000 6 Do[51]
port 95 nsew signal output
rlabel metal2 s 142784 159200 142840 160000 6 Do[52]
port 96 nsew signal output
rlabel metal2 s 144256 159200 144312 160000 6 Do[53]
port 97 nsew signal output
rlabel metal2 s 145636 159200 145692 160000 6 Do[54]
port 98 nsew signal output
rlabel metal2 s 147108 159200 147164 160000 6 Do[55]
port 99 nsew signal output
rlabel metal2 s 148488 159200 148544 160000 6 Do[56]
port 100 nsew signal output
rlabel metal2 s 149960 159200 150016 160000 6 Do[57]
port 101 nsew signal output
rlabel metal2 s 151340 159200 151396 160000 6 Do[58]
port 102 nsew signal output
rlabel metal2 s 152812 159200 152868 160000 6 Do[59]
port 103 nsew signal output
rlabel metal2 s 75624 159200 75680 160000 6 Do[5]
port 104 nsew signal output
rlabel metal2 s 154192 159200 154248 160000 6 Do[60]
port 105 nsew signal output
rlabel metal2 s 155664 159200 155720 160000 6 Do[61]
port 106 nsew signal output
rlabel metal2 s 157044 159200 157100 160000 6 Do[62]
port 107 nsew signal output
rlabel metal2 s 158516 159200 158572 160000 6 Do[63]
port 108 nsew signal output
rlabel metal2 s 77096 159200 77152 160000 6 Do[6]
port 109 nsew signal output
rlabel metal2 s 78476 159200 78532 160000 6 Do[7]
port 110 nsew signal output
rlabel metal2 s 79948 159200 80004 160000 6 Do[8]
port 111 nsew signal output
rlabel metal2 s 81420 159200 81476 160000 6 Do[9]
port 112 nsew signal output
rlabel metal2 s 19320 0 19376 800 6 clk
port 113 nsew signal input
rlabel metal2 s 139288 0 139344 800 6 hit
port 114 nsew signal output
rlabel metal3 s 158538 552 159338 672 6 line[0]
port 115 nsew signal input
rlabel metal3 s 158538 125400 159338 125520 6 line[100]
port 116 nsew signal input
rlabel metal3 s 158538 126624 159338 126744 6 line[101]
port 117 nsew signal input
rlabel metal3 s 158538 127984 159338 128104 6 line[102]
port 118 nsew signal input
rlabel metal3 s 158538 129208 159338 129328 6 line[103]
port 119 nsew signal input
rlabel metal3 s 158538 130432 159338 130552 6 line[104]
port 120 nsew signal input
rlabel metal3 s 158538 131656 159338 131776 6 line[105]
port 121 nsew signal input
rlabel metal3 s 158538 132880 159338 133000 6 line[106]
port 122 nsew signal input
rlabel metal3 s 158538 134240 159338 134360 6 line[107]
port 123 nsew signal input
rlabel metal3 s 158538 135464 159338 135584 6 line[108]
port 124 nsew signal input
rlabel metal3 s 158538 136688 159338 136808 6 line[109]
port 125 nsew signal input
rlabel metal3 s 158538 12928 159338 13048 6 line[10]
port 126 nsew signal input
rlabel metal3 s 158538 137912 159338 138032 6 line[110]
port 127 nsew signal input
rlabel metal3 s 158538 139136 159338 139256 6 line[111]
port 128 nsew signal input
rlabel metal3 s 158538 140496 159338 140616 6 line[112]
port 129 nsew signal input
rlabel metal3 s 158538 141720 159338 141840 6 line[113]
port 130 nsew signal input
rlabel metal3 s 158538 142944 159338 143064 6 line[114]
port 131 nsew signal input
rlabel metal3 s 158538 144168 159338 144288 6 line[115]
port 132 nsew signal input
rlabel metal3 s 158538 145392 159338 145512 6 line[116]
port 133 nsew signal input
rlabel metal3 s 158538 146616 159338 146736 6 line[117]
port 134 nsew signal input
rlabel metal3 s 158538 147976 159338 148096 6 line[118]
port 135 nsew signal input
rlabel metal3 s 158538 149200 159338 149320 6 line[119]
port 136 nsew signal input
rlabel metal3 s 158538 14288 159338 14408 6 line[11]
port 137 nsew signal input
rlabel metal3 s 158538 150424 159338 150544 6 line[120]
port 138 nsew signal input
rlabel metal3 s 158538 151648 159338 151768 6 line[121]
port 139 nsew signal input
rlabel metal3 s 158538 152872 159338 152992 6 line[122]
port 140 nsew signal input
rlabel metal3 s 158538 154232 159338 154352 6 line[123]
port 141 nsew signal input
rlabel metal3 s 158538 155456 159338 155576 6 line[124]
port 142 nsew signal input
rlabel metal3 s 158538 156680 159338 156800 6 line[125]
port 143 nsew signal input
rlabel metal3 s 158538 157904 159338 158024 6 line[126]
port 144 nsew signal input
rlabel metal3 s 158538 159128 159338 159248 6 line[127]
port 145 nsew signal input
rlabel metal3 s 158538 15512 159338 15632 6 line[12]
port 146 nsew signal input
rlabel metal3 s 158538 16736 159338 16856 6 line[13]
port 147 nsew signal input
rlabel metal3 s 158538 17960 159338 18080 6 line[14]
port 148 nsew signal input
rlabel metal3 s 158538 19184 159338 19304 6 line[15]
port 149 nsew signal input
rlabel metal3 s 158538 20544 159338 20664 6 line[16]
port 150 nsew signal input
rlabel metal3 s 158538 21768 159338 21888 6 line[17]
port 151 nsew signal input
rlabel metal3 s 158538 22992 159338 23112 6 line[18]
port 152 nsew signal input
rlabel metal3 s 158538 24216 159338 24336 6 line[19]
port 153 nsew signal input
rlabel metal3 s 158538 1776 159338 1896 6 line[1]
port 154 nsew signal input
rlabel metal3 s 158538 25440 159338 25560 6 line[20]
port 155 nsew signal input
rlabel metal3 s 158538 26664 159338 26784 6 line[21]
port 156 nsew signal input
rlabel metal3 s 158538 28024 159338 28144 6 line[22]
port 157 nsew signal input
rlabel metal3 s 158538 29248 159338 29368 6 line[23]
port 158 nsew signal input
rlabel metal3 s 158538 30472 159338 30592 6 line[24]
port 159 nsew signal input
rlabel metal3 s 158538 31696 159338 31816 6 line[25]
port 160 nsew signal input
rlabel metal3 s 158538 32920 159338 33040 6 line[26]
port 161 nsew signal input
rlabel metal3 s 158538 34280 159338 34400 6 line[27]
port 162 nsew signal input
rlabel metal3 s 158538 35504 159338 35624 6 line[28]
port 163 nsew signal input
rlabel metal3 s 158538 36728 159338 36848 6 line[29]
port 164 nsew signal input
rlabel metal3 s 158538 3000 159338 3120 6 line[2]
port 165 nsew signal input
rlabel metal3 s 158538 37952 159338 38072 6 line[30]
port 166 nsew signal input
rlabel metal3 s 158538 39176 159338 39296 6 line[31]
port 167 nsew signal input
rlabel metal3 s 158538 40536 159338 40656 6 line[32]
port 168 nsew signal input
rlabel metal3 s 158538 41760 159338 41880 6 line[33]
port 169 nsew signal input
rlabel metal3 s 158538 42984 159338 43104 6 line[34]
port 170 nsew signal input
rlabel metal3 s 158538 44208 159338 44328 6 line[35]
port 171 nsew signal input
rlabel metal3 s 158538 45432 159338 45552 6 line[36]
port 172 nsew signal input
rlabel metal3 s 158538 46656 159338 46776 6 line[37]
port 173 nsew signal input
rlabel metal3 s 158538 48016 159338 48136 6 line[38]
port 174 nsew signal input
rlabel metal3 s 158538 49240 159338 49360 6 line[39]
port 175 nsew signal input
rlabel metal3 s 158538 4224 159338 4344 6 line[3]
port 176 nsew signal input
rlabel metal3 s 158538 50464 159338 50584 6 line[40]
port 177 nsew signal input
rlabel metal3 s 158538 51688 159338 51808 6 line[41]
port 178 nsew signal input
rlabel metal3 s 158538 52912 159338 53032 6 line[42]
port 179 nsew signal input
rlabel metal3 s 158538 54272 159338 54392 6 line[43]
port 180 nsew signal input
rlabel metal3 s 158538 55496 159338 55616 6 line[44]
port 181 nsew signal input
rlabel metal3 s 158538 56720 159338 56840 6 line[45]
port 182 nsew signal input
rlabel metal3 s 158538 57944 159338 58064 6 line[46]
port 183 nsew signal input
rlabel metal3 s 158538 59168 159338 59288 6 line[47]
port 184 nsew signal input
rlabel metal3 s 158538 60528 159338 60648 6 line[48]
port 185 nsew signal input
rlabel metal3 s 158538 61752 159338 61872 6 line[49]
port 186 nsew signal input
rlabel metal3 s 158538 5448 159338 5568 6 line[4]
port 187 nsew signal input
rlabel metal3 s 158538 62976 159338 63096 6 line[50]
port 188 nsew signal input
rlabel metal3 s 158538 64200 159338 64320 6 line[51]
port 189 nsew signal input
rlabel metal3 s 158538 65424 159338 65544 6 line[52]
port 190 nsew signal input
rlabel metal3 s 158538 66648 159338 66768 6 line[53]
port 191 nsew signal input
rlabel metal3 s 158538 68008 159338 68128 6 line[54]
port 192 nsew signal input
rlabel metal3 s 158538 69232 159338 69352 6 line[55]
port 193 nsew signal input
rlabel metal3 s 158538 70456 159338 70576 6 line[56]
port 194 nsew signal input
rlabel metal3 s 158538 71680 159338 71800 6 line[57]
port 195 nsew signal input
rlabel metal3 s 158538 72904 159338 73024 6 line[58]
port 196 nsew signal input
rlabel metal3 s 158538 74264 159338 74384 6 line[59]
port 197 nsew signal input
rlabel metal3 s 158538 6672 159338 6792 6 line[5]
port 198 nsew signal input
rlabel metal3 s 158538 75488 159338 75608 6 line[60]
port 199 nsew signal input
rlabel metal3 s 158538 76712 159338 76832 6 line[61]
port 200 nsew signal input
rlabel metal3 s 158538 77936 159338 78056 6 line[62]
port 201 nsew signal input
rlabel metal3 s 158538 79160 159338 79280 6 line[63]
port 202 nsew signal input
rlabel metal3 s 158538 80520 159338 80640 6 line[64]
port 203 nsew signal input
rlabel metal3 s 158538 81744 159338 81864 6 line[65]
port 204 nsew signal input
rlabel metal3 s 158538 82968 159338 83088 6 line[66]
port 205 nsew signal input
rlabel metal3 s 158538 84192 159338 84312 6 line[67]
port 206 nsew signal input
rlabel metal3 s 158538 85416 159338 85536 6 line[68]
port 207 nsew signal input
rlabel metal3 s 158538 86640 159338 86760 6 line[69]
port 208 nsew signal input
rlabel metal3 s 158538 8032 159338 8152 6 line[6]
port 209 nsew signal input
rlabel metal3 s 158538 88000 159338 88120 6 line[70]
port 210 nsew signal input
rlabel metal3 s 158538 89224 159338 89344 6 line[71]
port 211 nsew signal input
rlabel metal3 s 158538 90448 159338 90568 6 line[72]
port 212 nsew signal input
rlabel metal3 s 158538 91672 159338 91792 6 line[73]
port 213 nsew signal input
rlabel metal3 s 158538 92896 159338 93016 6 line[74]
port 214 nsew signal input
rlabel metal3 s 158538 94256 159338 94376 6 line[75]
port 215 nsew signal input
rlabel metal3 s 158538 95480 159338 95600 6 line[76]
port 216 nsew signal input
rlabel metal3 s 158538 96704 159338 96824 6 line[77]
port 217 nsew signal input
rlabel metal3 s 158538 97928 159338 98048 6 line[78]
port 218 nsew signal input
rlabel metal3 s 158538 99152 159338 99272 6 line[79]
port 219 nsew signal input
rlabel metal3 s 158538 9256 159338 9376 6 line[7]
port 220 nsew signal input
rlabel metal3 s 158538 100512 159338 100632 6 line[80]
port 221 nsew signal input
rlabel metal3 s 158538 101736 159338 101856 6 line[81]
port 222 nsew signal input
rlabel metal3 s 158538 102960 159338 103080 6 line[82]
port 223 nsew signal input
rlabel metal3 s 158538 104184 159338 104304 6 line[83]
port 224 nsew signal input
rlabel metal3 s 158538 105408 159338 105528 6 line[84]
port 225 nsew signal input
rlabel metal3 s 158538 106632 159338 106752 6 line[85]
port 226 nsew signal input
rlabel metal3 s 158538 107992 159338 108112 6 line[86]
port 227 nsew signal input
rlabel metal3 s 158538 109216 159338 109336 6 line[87]
port 228 nsew signal input
rlabel metal3 s 158538 110440 159338 110560 6 line[88]
port 229 nsew signal input
rlabel metal3 s 158538 111664 159338 111784 6 line[89]
port 230 nsew signal input
rlabel metal3 s 158538 10480 159338 10600 6 line[8]
port 231 nsew signal input
rlabel metal3 s 158538 112888 159338 113008 6 line[90]
port 232 nsew signal input
rlabel metal3 s 158538 114248 159338 114368 6 line[91]
port 233 nsew signal input
rlabel metal3 s 158538 115472 159338 115592 6 line[92]
port 234 nsew signal input
rlabel metal3 s 158538 116696 159338 116816 6 line[93]
port 235 nsew signal input
rlabel metal3 s 158538 117920 159338 118040 6 line[94]
port 236 nsew signal input
rlabel metal3 s 158538 119144 159338 119264 6 line[95]
port 237 nsew signal input
rlabel metal3 s 158538 120504 159338 120624 6 line[96]
port 238 nsew signal input
rlabel metal3 s 158538 121728 159338 121848 6 line[97]
port 239 nsew signal input
rlabel metal3 s 158538 122952 159338 123072 6 line[98]
port 240 nsew signal input
rlabel metal3 s 158538 124176 159338 124296 6 line[99]
port 241 nsew signal input
rlabel metal3 s 158538 11704 159338 11824 6 line[9]
port 242 nsew signal input
rlabel metal2 s 59248 0 59304 800 6 rst_n
port 243 nsew signal input
rlabel metal2 s 99268 0 99324 800 6 wr
port 244 nsew signal input
rlabel metal4 s 157146 2128 157466 157808 6 VPWR
port 245 nsew power bidirectional
rlabel metal4 s 126426 2128 126746 157808 6 VPWR
port 246 nsew power bidirectional
rlabel metal4 s 95706 2128 96026 157808 6 VPWR
port 247 nsew power bidirectional
rlabel metal4 s 64986 2128 65306 157808 6 VPWR
port 248 nsew power bidirectional
rlabel metal4 s 34266 2128 34586 157808 6 VPWR
port 249 nsew power bidirectional
rlabel metal4 s 3546 2128 3866 157808 6 VPWR
port 250 nsew power bidirectional
rlabel metal4 s 141786 2128 142106 157808 6 VGND
port 251 nsew ground bidirectional
rlabel metal4 s 111066 2128 111386 157808 6 VGND
port 252 nsew ground bidirectional
rlabel metal4 s 80346 2128 80666 157808 6 VGND
port 253 nsew ground bidirectional
rlabel metal4 s 49626 2128 49946 157808 6 VGND
port 254 nsew ground bidirectional
rlabel metal4 s 18906 2128 19226 157808 6 VGND
port 255 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 159338 160000
string LEFview TRUE
<< end >>
